magic
tech sky130B
magscale 1 2
timestamp 1662560833
<< viali >>
rect 4905 47141 4939 47175
rect 27813 47141 27847 47175
rect 47041 47141 47075 47175
rect 1409 47073 1443 47107
rect 1685 47005 1719 47039
rect 2789 47005 2823 47039
rect 4261 47005 4295 47039
rect 5549 47005 5583 47039
rect 9137 47005 9171 47039
rect 12725 47005 12759 47039
rect 13461 47005 13495 47039
rect 14473 47005 14507 47039
rect 15669 47005 15703 47039
rect 24869 47005 24903 47039
rect 25513 47005 25547 47039
rect 26433 47005 26467 47039
rect 27997 47005 28031 47039
rect 30113 47005 30147 47039
rect 33057 47005 33091 47039
rect 36093 47005 36127 47039
rect 46397 47005 46431 47039
rect 47593 47005 47627 47039
rect 2881 46937 2915 46971
rect 47685 46937 47719 46971
rect 8953 46869 8987 46903
rect 1869 46597 1903 46631
rect 3985 46529 4019 46563
rect 11897 46529 11931 46563
rect 14197 46529 14231 46563
rect 24593 46529 24627 46563
rect 26985 46529 27019 46563
rect 29745 46529 29779 46563
rect 32781 46529 32815 46563
rect 35817 46529 35851 46563
rect 37289 46529 37323 46563
rect 45201 46529 45235 46563
rect 47593 46529 47627 46563
rect 1685 46461 1719 46495
rect 2145 46461 2179 46495
rect 4169 46461 4203 46495
rect 4629 46461 4663 46495
rect 12081 46461 12115 46495
rect 12909 46461 12943 46495
rect 14381 46461 14415 46495
rect 14841 46461 14875 46495
rect 22293 46461 22327 46495
rect 22477 46461 22511 46495
rect 23213 46461 23247 46495
rect 24777 46461 24811 46495
rect 25789 46461 25823 46495
rect 27169 46461 27203 46495
rect 27629 46461 27663 46495
rect 29929 46461 29963 46495
rect 30389 46461 30423 46495
rect 32965 46461 32999 46495
rect 33517 46461 33551 46495
rect 37473 46461 37507 46495
rect 37749 46461 37783 46495
rect 45385 46461 45419 46495
rect 46765 46461 46799 46495
rect 36645 46393 36679 46427
rect 10977 46325 11011 46359
rect 35909 46325 35943 46359
rect 41797 46325 41831 46359
rect 47685 46325 47719 46359
rect 4169 46121 4203 46155
rect 14473 46121 14507 46155
rect 23029 46121 23063 46155
rect 32873 46121 32907 46155
rect 2789 45985 2823 46019
rect 5273 45985 5307 46019
rect 5825 45985 5859 46019
rect 9597 45985 9631 46019
rect 10885 45985 10919 46019
rect 11345 45985 11379 46019
rect 15393 45985 15427 46019
rect 15853 45985 15887 46019
rect 36185 45985 36219 46019
rect 41613 45985 41647 46019
rect 42073 45985 42107 46019
rect 48145 45985 48179 46019
rect 1409 45917 1443 45951
rect 4077 45917 4111 45951
rect 9229 45917 9263 45951
rect 13185 45917 13219 45951
rect 14381 45917 14415 45951
rect 24685 45917 24719 45951
rect 26985 45917 27019 45951
rect 28825 45917 28859 45951
rect 29745 45917 29779 45951
rect 32781 45917 32815 45951
rect 35725 45917 35759 45951
rect 38301 45917 38335 45951
rect 45845 45917 45879 45951
rect 46305 45917 46339 45951
rect 1593 45849 1627 45883
rect 5457 45849 5491 45883
rect 11069 45849 11103 45883
rect 15577 45849 15611 45883
rect 24869 45849 24903 45883
rect 26525 45849 26559 45883
rect 27169 45849 27203 45883
rect 35909 45849 35943 45883
rect 41797 45849 41831 45883
rect 46489 45849 46523 45883
rect 13277 45781 13311 45815
rect 11621 45577 11655 45611
rect 15669 45577 15703 45611
rect 22937 45577 22971 45611
rect 1685 45509 1719 45543
rect 2513 45509 2547 45543
rect 5549 45509 5583 45543
rect 12633 45509 12667 45543
rect 13369 45509 13403 45543
rect 24685 45509 24719 45543
rect 25329 45509 25363 45543
rect 39957 45509 39991 45543
rect 45385 45509 45419 45543
rect 47685 45509 47719 45543
rect 5457 45441 5491 45475
rect 8401 45441 8435 45475
rect 8585 45441 8619 45475
rect 9137 45441 9171 45475
rect 10333 45441 10367 45475
rect 11529 45441 11563 45475
rect 12541 45441 12575 45475
rect 13185 45441 13219 45475
rect 15577 45441 15611 45475
rect 22845 45441 22879 45475
rect 24593 45441 24627 45475
rect 25237 45441 25271 45475
rect 26065 45441 26099 45475
rect 26157 45441 26191 45475
rect 27261 45441 27295 45475
rect 28641 45441 28675 45475
rect 35933 45441 35967 45475
rect 38117 45441 38151 45475
rect 45201 45441 45235 45475
rect 47593 45441 47627 45475
rect 2329 45373 2363 45407
rect 3065 45373 3099 45407
rect 9413 45373 9447 45407
rect 10885 45373 10919 45407
rect 14289 45373 14323 45407
rect 28825 45373 28859 45407
rect 30297 45373 30331 45407
rect 38301 45373 38335 45407
rect 46857 45373 46891 45407
rect 1869 45305 1903 45339
rect 36001 45305 36035 45339
rect 1961 45033 1995 45067
rect 3157 45033 3191 45067
rect 3893 45033 3927 45067
rect 26801 45033 26835 45067
rect 27445 45033 27479 45067
rect 30021 45033 30055 45067
rect 38209 45033 38243 45067
rect 41797 45033 41831 45067
rect 2605 44965 2639 44999
rect 48145 44897 48179 44931
rect 3065 44829 3099 44863
rect 3801 44829 3835 44863
rect 9229 44829 9263 44863
rect 26709 44829 26743 44863
rect 27353 44829 27387 44863
rect 29929 44829 29963 44863
rect 38117 44829 38151 44863
rect 41705 44829 41739 44863
rect 45845 44829 45879 44863
rect 46305 44829 46339 44863
rect 9597 44761 9631 44795
rect 46489 44761 46523 44795
rect 46305 44489 46339 44523
rect 9137 44353 9171 44387
rect 46213 44353 46247 44387
rect 47593 44353 47627 44387
rect 9413 44285 9447 44319
rect 47685 44217 47719 44251
rect 47041 44149 47075 44183
rect 48053 43809 48087 43843
rect 2329 43741 2363 43775
rect 40417 43741 40451 43775
rect 46305 43741 46339 43775
rect 46489 43673 46523 43707
rect 46581 43401 46615 43435
rect 3985 43333 4019 43367
rect 2145 43265 2179 43299
rect 40049 43265 40083 43299
rect 46029 43265 46063 43299
rect 46489 43265 46523 43299
rect 47593 43265 47627 43299
rect 2329 43197 2363 43231
rect 40233 43197 40267 43231
rect 41429 43197 41463 43231
rect 47685 43061 47719 43095
rect 3893 42721 3927 42755
rect 26985 42721 27019 42755
rect 27997 42721 28031 42755
rect 46489 42721 46523 42755
rect 3801 42653 3835 42687
rect 27169 42653 27203 42687
rect 28181 42653 28215 42687
rect 33701 42653 33735 42687
rect 45201 42653 45235 42687
rect 45845 42653 45879 42687
rect 46305 42653 46339 42687
rect 27721 42585 27755 42619
rect 48145 42585 48179 42619
rect 27353 42517 27387 42551
rect 28365 42517 28399 42551
rect 33517 42517 33551 42551
rect 45017 42517 45051 42551
rect 40325 42313 40359 42347
rect 33416 42245 33450 42279
rect 37657 42245 37691 42279
rect 45385 42245 45419 42279
rect 27169 42177 27203 42211
rect 28549 42177 28583 42211
rect 31401 42177 31435 42211
rect 32689 42177 32723 42211
rect 35173 42177 35207 42211
rect 35357 42177 35391 42211
rect 36001 42177 36035 42211
rect 36645 42177 36679 42211
rect 37473 42177 37507 42211
rect 40233 42177 40267 42211
rect 41613 42177 41647 42211
rect 41705 42177 41739 42211
rect 42533 42177 42567 42211
rect 42625 42177 42659 42211
rect 42809 42177 42843 42211
rect 43453 42177 43487 42211
rect 45201 42177 45235 42211
rect 33149 42109 33183 42143
rect 34989 42109 35023 42143
rect 37289 42109 37323 42143
rect 46857 42109 46891 42143
rect 26985 41973 27019 42007
rect 28365 41973 28399 42007
rect 31217 41973 31251 42007
rect 32505 41973 32539 42007
rect 34529 41973 34563 42007
rect 35817 41973 35851 42007
rect 36461 41973 36495 42007
rect 41889 41973 41923 42007
rect 43269 41973 43303 42007
rect 47777 41973 47811 42007
rect 33609 41769 33643 41803
rect 36645 41769 36679 41803
rect 42533 41769 42567 41803
rect 35265 41633 35299 41667
rect 46305 41633 46339 41667
rect 26525 41565 26559 41599
rect 29561 41565 29595 41599
rect 29817 41565 29851 41599
rect 31401 41565 31435 41599
rect 33333 41565 33367 41599
rect 33425 41565 33459 41599
rect 35532 41565 35566 41599
rect 37105 41565 37139 41599
rect 39313 41565 39347 41599
rect 39865 41565 39899 41599
rect 40049 41565 40083 41599
rect 41153 41565 41187 41599
rect 42993 41565 43027 41599
rect 45109 41565 45143 41599
rect 45293 41565 45327 41599
rect 26792 41497 26826 41531
rect 31646 41497 31680 41531
rect 37350 41497 37384 41531
rect 40233 41497 40267 41531
rect 41420 41497 41454 41531
rect 43260 41497 43294 41531
rect 46489 41497 46523 41531
rect 48145 41497 48179 41531
rect 27905 41429 27939 41463
rect 30941 41429 30975 41463
rect 32781 41429 32815 41463
rect 38485 41429 38519 41463
rect 39129 41429 39163 41463
rect 44373 41429 44407 41463
rect 45477 41429 45511 41463
rect 31217 41225 31251 41259
rect 34437 41225 34471 41259
rect 39405 41225 39439 41259
rect 41705 41225 41739 41259
rect 42717 41225 42751 41259
rect 45385 41225 45419 41259
rect 46949 41225 46983 41259
rect 9045 41157 9079 41191
rect 17049 41157 17083 41191
rect 32658 41157 32692 41191
rect 34529 41157 34563 41191
rect 36277 41157 36311 41191
rect 40132 41157 40166 41191
rect 42441 41157 42475 41191
rect 16957 41089 16991 41123
rect 25513 41089 25547 41123
rect 26157 41089 26191 41123
rect 29561 41089 29595 41123
rect 31033 41089 31067 41123
rect 34621 41089 34655 41123
rect 35265 41089 35299 41123
rect 35541 41089 35575 41123
rect 36553 41089 36587 41123
rect 37565 41089 37599 41123
rect 38025 41089 38059 41123
rect 38281 41089 38315 41123
rect 41889 41089 41923 41123
rect 42625 41089 42659 41123
rect 42809 41089 42843 41123
rect 44005 41089 44039 41123
rect 44261 41089 44295 41123
rect 46029 41089 46063 41123
rect 46857 41089 46891 41123
rect 8861 41021 8895 41055
rect 9321 41021 9355 41055
rect 25973 41021 26007 41055
rect 30849 41021 30883 41055
rect 32413 41021 32447 41055
rect 35357 41021 35391 41055
rect 36461 41021 36495 41055
rect 39865 41021 39899 41055
rect 26341 40953 26375 40987
rect 33793 40953 33827 40987
rect 34253 40953 34287 40987
rect 37381 40953 37415 40987
rect 25329 40885 25363 40919
rect 29377 40885 29411 40919
rect 34805 40885 34839 40919
rect 35265 40885 35299 40919
rect 35725 40885 35759 40919
rect 36553 40885 36587 40919
rect 36737 40885 36771 40919
rect 41245 40885 41279 40919
rect 42993 40885 43027 40919
rect 45845 40885 45879 40919
rect 47777 40885 47811 40919
rect 9137 40681 9171 40715
rect 27905 40681 27939 40715
rect 29009 40681 29043 40715
rect 33793 40681 33827 40715
rect 38393 40681 38427 40715
rect 38853 40681 38887 40715
rect 41613 40681 41647 40715
rect 42073 40681 42107 40715
rect 22753 40545 22787 40579
rect 28641 40545 28675 40579
rect 29561 40545 29595 40579
rect 42257 40545 42291 40579
rect 42993 40545 43027 40579
rect 46305 40545 46339 40579
rect 23213 40477 23247 40511
rect 23305 40477 23339 40511
rect 24593 40477 24627 40511
rect 25053 40477 25087 40511
rect 25320 40477 25354 40511
rect 26985 40477 27019 40511
rect 27077 40477 27111 40511
rect 27905 40477 27939 40511
rect 27997 40477 28031 40511
rect 28825 40477 28859 40511
rect 29817 40477 29851 40511
rect 33517 40477 33551 40511
rect 33609 40477 33643 40511
rect 34989 40477 35023 40511
rect 35173 40477 35207 40511
rect 36553 40477 36587 40511
rect 37013 40477 37047 40511
rect 38117 40477 38151 40511
rect 38209 40477 38243 40511
rect 39037 40477 39071 40511
rect 40233 40477 40267 40511
rect 42349 40477 42383 40511
rect 43177 40477 43211 40511
rect 43821 40477 43855 40511
rect 44005 40477 44039 40511
rect 27721 40409 27755 40443
rect 37381 40409 37415 40443
rect 37565 40409 37599 40443
rect 40500 40409 40534 40443
rect 42073 40409 42107 40443
rect 46489 40409 46523 40443
rect 48145 40409 48179 40443
rect 23489 40341 23523 40375
rect 24409 40341 24443 40375
rect 26433 40341 26467 40375
rect 27261 40341 27295 40375
rect 28181 40341 28215 40375
rect 30941 40341 30975 40375
rect 35357 40341 35391 40375
rect 36369 40341 36403 40375
rect 37197 40341 37231 40375
rect 37289 40341 37323 40375
rect 42533 40341 42567 40375
rect 43361 40341 43395 40375
rect 44189 40341 44223 40375
rect 25881 40137 25915 40171
rect 43913 40137 43947 40171
rect 46397 40137 46431 40171
rect 24746 40069 24780 40103
rect 23857 40001 23891 40035
rect 27169 40001 27203 40035
rect 27436 40001 27470 40035
rect 29193 40001 29227 40035
rect 30205 40001 30239 40035
rect 44097 40001 44131 40035
rect 45284 40001 45318 40035
rect 46857 40001 46891 40035
rect 46949 40001 46983 40035
rect 24501 39933 24535 39967
rect 45017 39933 45051 39967
rect 29009 39865 29043 39899
rect 23673 39797 23707 39831
rect 28549 39797 28583 39831
rect 30021 39797 30055 39831
rect 47777 39797 47811 39831
rect 26617 39593 26651 39627
rect 28641 39593 28675 39627
rect 32597 39593 32631 39627
rect 27629 39525 27663 39559
rect 26249 39457 26283 39491
rect 46305 39457 46339 39491
rect 24409 39389 24443 39423
rect 26433 39389 26467 39423
rect 27905 39389 27939 39423
rect 28825 39389 28859 39423
rect 30757 39389 30791 39423
rect 30849 39389 30883 39423
rect 31033 39389 31067 39423
rect 31677 39389 31711 39423
rect 32413 39389 32447 39423
rect 34989 39389 35023 39423
rect 35081 39389 35115 39423
rect 35311 39389 35345 39423
rect 35449 39389 35483 39423
rect 41889 39389 41923 39423
rect 42993 39389 43027 39423
rect 24654 39321 24688 39355
rect 27997 39321 28031 39355
rect 35173 39321 35207 39355
rect 41705 39321 41739 39355
rect 46489 39321 46523 39355
rect 48145 39321 48179 39355
rect 25789 39253 25823 39287
rect 27813 39253 27847 39287
rect 28181 39253 28215 39287
rect 31493 39253 31527 39287
rect 34805 39253 34839 39287
rect 42073 39253 42107 39287
rect 42809 39253 42843 39287
rect 36369 39049 36403 39083
rect 41061 39049 41095 39083
rect 41153 39049 41187 39083
rect 47685 39049 47719 39083
rect 33968 38981 34002 39015
rect 39221 38981 39255 39015
rect 39451 38981 39485 39015
rect 40969 38981 41003 39015
rect 30021 38913 30055 38947
rect 32321 38913 32355 38947
rect 35725 38913 35759 38947
rect 35909 38913 35943 38947
rect 36553 38913 36587 38947
rect 37565 38913 37599 38947
rect 37749 38913 37783 38947
rect 38393 38913 38427 38947
rect 39129 38913 39163 38947
rect 39313 38913 39347 38947
rect 40233 38913 40267 38947
rect 42441 38913 42475 38947
rect 42708 38913 42742 38947
rect 45201 38913 45235 38947
rect 45468 38913 45502 38947
rect 47593 38913 47627 38947
rect 29837 38845 29871 38879
rect 30757 38845 30791 38879
rect 31033 38845 31067 38879
rect 32137 38845 32171 38879
rect 33701 38845 33735 38879
rect 35541 38845 35575 38879
rect 37381 38845 37415 38879
rect 39589 38845 39623 38879
rect 41337 38845 41371 38879
rect 38209 38777 38243 38811
rect 40785 38777 40819 38811
rect 30205 38709 30239 38743
rect 32505 38709 32539 38743
rect 35081 38709 35115 38743
rect 38945 38709 38979 38743
rect 40049 38709 40083 38743
rect 43821 38709 43855 38743
rect 46581 38709 46615 38743
rect 42073 38505 42107 38539
rect 42349 38505 42383 38539
rect 46765 38505 46799 38539
rect 32229 38437 32263 38471
rect 30389 38369 30423 38403
rect 34713 38369 34747 38403
rect 42073 38369 42107 38403
rect 45937 38369 45971 38403
rect 25789 38301 25823 38335
rect 28733 38301 28767 38335
rect 30021 38301 30055 38335
rect 30849 38301 30883 38335
rect 32873 38301 32907 38335
rect 34969 38301 35003 38335
rect 37197 38301 37231 38335
rect 37464 38301 37498 38335
rect 40049 38301 40083 38335
rect 42165 38301 42199 38335
rect 43085 38301 43119 38335
rect 45109 38301 45143 38335
rect 45201 38301 45235 38335
rect 46121 38301 46155 38335
rect 46949 38301 46983 38335
rect 47409 38301 47443 38335
rect 28549 38233 28583 38267
rect 29837 38233 29871 38267
rect 31116 38233 31150 38267
rect 40316 38233 40350 38267
rect 41889 38233 41923 38267
rect 43352 38233 43386 38267
rect 45385 38233 45419 38267
rect 25605 38165 25639 38199
rect 28917 38165 28951 38199
rect 30113 38165 30147 38199
rect 30205 38165 30239 38199
rect 32689 38165 32723 38199
rect 36093 38165 36127 38199
rect 38577 38165 38611 38199
rect 41429 38165 41463 38199
rect 44465 38165 44499 38199
rect 46305 38165 46339 38199
rect 47501 38165 47535 38199
rect 30573 37961 30607 37995
rect 35633 37961 35667 37995
rect 38669 37961 38703 37995
rect 40969 37961 41003 37995
rect 41797 37961 41831 37995
rect 43913 37961 43947 37995
rect 47593 37961 47627 37995
rect 32404 37893 32438 37927
rect 35842 37893 35876 37927
rect 45928 37893 45962 37927
rect 25320 37825 25354 37859
rect 29193 37825 29227 37859
rect 29460 37825 29494 37859
rect 31033 37825 31067 37859
rect 31217 37825 31251 37859
rect 31309 37825 31343 37859
rect 35725 37825 35759 37859
rect 36461 37825 36495 37859
rect 36645 37825 36679 37859
rect 37289 37825 37323 37859
rect 37556 37825 37590 37859
rect 39856 37825 39890 37859
rect 41429 37825 41463 37859
rect 41613 37825 41647 37859
rect 44097 37825 44131 37859
rect 45661 37825 45695 37859
rect 47777 37825 47811 37859
rect 25053 37757 25087 37791
rect 32137 37757 32171 37791
rect 35357 37757 35391 37791
rect 39589 37757 39623 37791
rect 31493 37689 31527 37723
rect 26433 37621 26467 37655
rect 31033 37621 31067 37655
rect 33517 37621 33551 37655
rect 36001 37621 36035 37655
rect 36461 37621 36495 37655
rect 47041 37621 47075 37655
rect 26157 37417 26191 37451
rect 29653 37417 29687 37451
rect 41521 37417 41555 37451
rect 35817 37349 35851 37383
rect 36737 37349 36771 37383
rect 26801 37281 26835 37315
rect 29009 37281 29043 37315
rect 34713 37281 34747 37315
rect 35541 37281 35575 37315
rect 39865 37281 39899 37315
rect 40693 37281 40727 37315
rect 24961 37213 24995 37247
rect 25789 37213 25823 37247
rect 25973 37213 26007 37247
rect 26985 37213 27019 37247
rect 27169 37213 27203 37247
rect 27813 37213 27847 37247
rect 28549 37213 28583 37247
rect 28641 37213 28675 37247
rect 28871 37213 28905 37247
rect 29837 37213 29871 37247
rect 34897 37213 34931 37247
rect 36461 37213 36495 37247
rect 40049 37213 40083 37247
rect 40877 37213 40911 37247
rect 41705 37213 41739 37247
rect 44005 37213 44039 37247
rect 44097 37213 44131 37247
rect 44281 37213 44315 37247
rect 46305 37213 46339 37247
rect 28733 37145 28767 37179
rect 40233 37145 40267 37179
rect 46489 37145 46523 37179
rect 48145 37145 48179 37179
rect 24777 37077 24811 37111
rect 27629 37077 27663 37111
rect 28365 37077 28399 37111
rect 35081 37077 35115 37111
rect 36001 37077 36035 37111
rect 36921 37077 36955 37111
rect 41061 37077 41095 37111
rect 36185 36873 36219 36907
rect 29070 36805 29104 36839
rect 44741 36805 44775 36839
rect 44957 36805 44991 36839
rect 24308 36737 24342 36771
rect 26985 36737 27019 36771
rect 27252 36737 27286 36771
rect 28825 36737 28859 36771
rect 33140 36737 33174 36771
rect 34989 36737 35023 36771
rect 35081 36737 35115 36771
rect 35265 36737 35299 36771
rect 35357 36737 35391 36771
rect 36001 36737 36035 36771
rect 36277 36737 36311 36771
rect 39037 36737 39071 36771
rect 41429 36737 41463 36771
rect 47041 36737 47075 36771
rect 47777 36737 47811 36771
rect 24041 36669 24075 36703
rect 32873 36669 32907 36703
rect 45109 36601 45143 36635
rect 25421 36533 25455 36567
rect 28365 36533 28399 36567
rect 30205 36533 30239 36567
rect 34253 36533 34287 36567
rect 34805 36533 34839 36567
rect 35817 36533 35851 36567
rect 40509 36533 40543 36567
rect 41245 36533 41279 36567
rect 44925 36533 44959 36567
rect 46857 36533 46891 36567
rect 25789 36329 25823 36363
rect 42257 36329 42291 36363
rect 46305 36329 46339 36363
rect 26801 36261 26835 36295
rect 40417 36261 40451 36295
rect 45753 36261 45787 36295
rect 29561 36193 29595 36227
rect 34713 36193 34747 36227
rect 36461 36193 36495 36227
rect 46765 36193 46799 36227
rect 19901 36125 19935 36159
rect 24409 36125 24443 36159
rect 24676 36125 24710 36159
rect 26985 36125 27019 36159
rect 27077 36125 27111 36159
rect 29745 36125 29779 36159
rect 34989 36125 35023 36159
rect 36185 36125 36219 36159
rect 36277 36125 36311 36159
rect 36553 36125 36587 36159
rect 40877 36125 40911 36159
rect 42717 36125 42751 36159
rect 45937 36125 45971 36159
rect 47021 36125 47055 36159
rect 20361 36057 20395 36091
rect 40233 36057 40267 36091
rect 41144 36057 41178 36091
rect 42984 36057 43018 36091
rect 46029 36057 46063 36091
rect 27169 35989 27203 36023
rect 27353 35989 27387 36023
rect 29929 35989 29963 36023
rect 36001 35989 36035 36023
rect 44097 35989 44131 36023
rect 46121 35989 46155 36023
rect 48145 35989 48179 36023
rect 24225 35785 24259 35819
rect 25237 35785 25271 35819
rect 39865 35785 39899 35819
rect 40693 35785 40727 35819
rect 42809 35785 42843 35819
rect 43913 35785 43947 35819
rect 46857 35785 46891 35819
rect 47961 35785 47995 35819
rect 25697 35717 25731 35751
rect 26985 35717 27019 35751
rect 39221 35717 39255 35751
rect 39681 35717 39715 35751
rect 44005 35717 44039 35751
rect 45477 35717 45511 35751
rect 24409 35649 24443 35683
rect 25053 35649 25087 35683
rect 25973 35649 26007 35683
rect 27261 35649 27295 35683
rect 29561 35649 29595 35683
rect 32321 35649 32355 35683
rect 35081 35649 35115 35683
rect 35265 35649 35299 35683
rect 35357 35649 35391 35683
rect 35449 35649 35483 35683
rect 35633 35649 35667 35683
rect 38945 35649 38979 35683
rect 39957 35649 39991 35683
rect 40877 35649 40911 35683
rect 42993 35649 43027 35683
rect 43637 35649 43671 35683
rect 44557 35649 44591 35683
rect 44741 35649 44775 35683
rect 44925 35649 44959 35683
rect 45753 35649 45787 35683
rect 46397 35649 46431 35683
rect 46673 35649 46707 35683
rect 47593 35649 47627 35683
rect 47777 35649 47811 35683
rect 24869 35581 24903 35615
rect 25789 35581 25823 35615
rect 27169 35581 27203 35615
rect 32413 35581 32447 35615
rect 39221 35581 39255 35615
rect 43729 35581 43763 35615
rect 44097 35581 44131 35615
rect 45017 35581 45051 35615
rect 45569 35581 45603 35615
rect 46581 35581 46615 35615
rect 45937 35513 45971 35547
rect 25973 35445 26007 35479
rect 26157 35445 26191 35479
rect 26985 35445 27019 35479
rect 27445 35445 27479 35479
rect 29377 35445 29411 35479
rect 32689 35445 32723 35479
rect 35817 35445 35851 35479
rect 39037 35445 39071 35479
rect 39681 35445 39715 35479
rect 43453 35445 43487 35479
rect 45477 35445 45511 35479
rect 46397 35445 46431 35479
rect 25237 35241 25271 35275
rect 44189 35241 44223 35275
rect 48145 35241 48179 35275
rect 35909 35173 35943 35207
rect 24869 35105 24903 35139
rect 38853 35105 38887 35139
rect 39313 35105 39347 35139
rect 43821 35105 43855 35139
rect 46765 35105 46799 35139
rect 2329 35037 2363 35071
rect 25053 35037 25087 35071
rect 26157 35037 26191 35071
rect 26249 35037 26283 35071
rect 26433 35037 26467 35071
rect 27721 35037 27755 35071
rect 27813 35037 27847 35071
rect 28181 35037 28215 35071
rect 30941 35037 30975 35071
rect 34713 35037 34747 35071
rect 34897 35037 34931 35071
rect 36185 35037 36219 35071
rect 36645 35037 36679 35071
rect 38945 35037 38979 35071
rect 39865 35037 39899 35071
rect 44005 35037 44039 35071
rect 45017 35037 45051 35071
rect 45201 35037 45235 35071
rect 46305 35037 46339 35071
rect 25881 34969 25915 35003
rect 27905 34969 27939 35003
rect 28023 34969 28057 35003
rect 31208 34969 31242 35003
rect 35909 34969 35943 35003
rect 36890 34969 36924 35003
rect 40132 34969 40166 35003
rect 47010 34969 47044 35003
rect 26065 34901 26099 34935
rect 27537 34901 27571 34935
rect 32321 34901 32355 34935
rect 34805 34901 34839 34935
rect 36093 34901 36127 34935
rect 38025 34901 38059 34935
rect 41245 34901 41279 34935
rect 45385 34901 45419 34935
rect 46121 34901 46155 34935
rect 25789 34697 25823 34731
rect 27445 34697 27479 34731
rect 32873 34697 32907 34731
rect 33517 34697 33551 34731
rect 37565 34697 37599 34731
rect 39405 34697 39439 34731
rect 45385 34697 45419 34731
rect 46857 34697 46891 34731
rect 27261 34629 27295 34663
rect 28150 34629 28184 34663
rect 29990 34629 30024 34663
rect 2053 34561 2087 34595
rect 24409 34561 24443 34595
rect 24665 34561 24699 34595
rect 27077 34561 27111 34595
rect 27905 34561 27939 34595
rect 32137 34561 32171 34595
rect 32321 34561 32355 34595
rect 32689 34561 32723 34595
rect 33425 34561 33459 34595
rect 33609 34561 33643 34595
rect 34253 34561 34287 34595
rect 34437 34561 34471 34595
rect 34529 34561 34563 34595
rect 34989 34561 35023 34595
rect 35173 34561 35207 34595
rect 35633 34561 35667 34595
rect 36553 34561 36587 34595
rect 37289 34561 37323 34595
rect 37381 34561 37415 34595
rect 39037 34561 39071 34595
rect 41153 34561 41187 34595
rect 44005 34561 44039 34595
rect 44272 34561 44306 34595
rect 46489 34561 46523 34595
rect 46673 34561 46707 34595
rect 2237 34493 2271 34527
rect 3617 34493 3651 34527
rect 29745 34493 29779 34527
rect 32413 34493 32447 34527
rect 32505 34493 32539 34527
rect 35725 34493 35759 34527
rect 36737 34493 36771 34527
rect 37565 34493 37599 34527
rect 39129 34493 39163 34527
rect 41245 34493 41279 34527
rect 29285 34357 29319 34391
rect 31125 34357 31159 34391
rect 34069 34357 34103 34391
rect 35081 34357 35115 34391
rect 2421 34153 2455 34187
rect 23673 34153 23707 34187
rect 27537 34153 27571 34187
rect 31309 34153 31343 34187
rect 33241 34153 33275 34187
rect 36645 34153 36679 34187
rect 41061 34153 41095 34187
rect 43821 34153 43855 34187
rect 45017 34153 45051 34187
rect 32137 34085 32171 34119
rect 24961 34017 24995 34051
rect 30757 34017 30791 34051
rect 32413 34017 32447 34051
rect 32505 34017 32539 34051
rect 36461 34017 36495 34051
rect 41705 34017 41739 34051
rect 43361 34017 43395 34051
rect 46765 34017 46799 34051
rect 2329 33949 2363 33983
rect 23857 33949 23891 33983
rect 24685 33949 24719 33983
rect 24777 33949 24811 33983
rect 29745 33949 29779 33983
rect 30665 33949 30699 33983
rect 30849 33949 30883 33983
rect 31585 33949 31619 33983
rect 32321 33949 32355 33983
rect 32597 33949 32631 33983
rect 33149 33949 33183 33983
rect 33333 33949 33367 33983
rect 33977 33949 34011 33983
rect 34713 33949 34747 33983
rect 36369 33949 36403 33983
rect 40693 33949 40727 33983
rect 40877 33949 40911 33983
rect 41521 33949 41555 33983
rect 44005 33949 44039 33983
rect 45201 33949 45235 33983
rect 26065 33881 26099 33915
rect 31309 33881 31343 33915
rect 31493 33881 31527 33915
rect 34161 33881 34195 33915
rect 34897 33881 34931 33915
rect 47032 33881 47066 33915
rect 29561 33813 29595 33847
rect 35081 33813 35115 33847
rect 48145 33813 48179 33847
rect 25513 33609 25547 33643
rect 25973 33609 26007 33643
rect 34713 33609 34747 33643
rect 41245 33609 41279 33643
rect 46857 33609 46891 33643
rect 30941 33541 30975 33575
rect 33241 33541 33275 33575
rect 34345 33541 34379 33575
rect 43076 33541 43110 33575
rect 24133 33473 24167 33507
rect 24400 33473 24434 33507
rect 26157 33473 26191 33507
rect 28641 33473 28675 33507
rect 31125 33473 31159 33507
rect 32413 33473 32447 33507
rect 32505 33473 32539 33507
rect 33517 33473 33551 33507
rect 33606 33473 33640 33507
rect 33701 33476 33735 33510
rect 33885 33473 33919 33507
rect 34529 33473 34563 33507
rect 34805 33473 34839 33507
rect 41429 33473 41463 33507
rect 42809 33473 42843 33507
rect 44833 33473 44867 33507
rect 47041 33473 47075 33507
rect 30297 33405 30331 33439
rect 32321 33405 32355 33439
rect 32597 33405 32631 33439
rect 44189 33337 44223 33371
rect 32137 33269 32171 33303
rect 44649 33269 44683 33303
rect 47777 33269 47811 33303
rect 24869 33065 24903 33099
rect 30389 33065 30423 33099
rect 31677 33065 31711 33099
rect 33057 33065 33091 33099
rect 37381 33065 37415 33099
rect 40049 33065 40083 33099
rect 40785 33065 40819 33099
rect 40969 33065 41003 33099
rect 42901 33065 42935 33099
rect 43821 33065 43855 33099
rect 47685 33065 47719 33099
rect 27629 32929 27663 32963
rect 30021 32929 30055 32963
rect 31401 32929 31435 32963
rect 35725 32929 35759 32963
rect 37105 32929 37139 32963
rect 45017 32929 45051 32963
rect 2329 32861 2363 32895
rect 24593 32861 24627 32895
rect 24685 32861 24719 32895
rect 25421 32861 25455 32895
rect 25513 32861 25547 32895
rect 26341 32861 26375 32895
rect 27896 32861 27930 32895
rect 30205 32861 30239 32895
rect 31309 32861 31343 32895
rect 32321 32861 32355 32895
rect 32597 32861 32631 32895
rect 33241 32861 33275 32895
rect 33425 32861 33459 32895
rect 33517 32861 33551 32895
rect 35541 32861 35575 32895
rect 37013 32861 37047 32895
rect 44005 32861 44039 32895
rect 45273 32861 45307 32895
rect 46857 32861 46891 32895
rect 47041 32861 47075 32895
rect 47225 32861 47259 32895
rect 47869 32861 47903 32895
rect 39957 32793 39991 32827
rect 40601 32793 40635 32827
rect 41613 32793 41647 32827
rect 25697 32725 25731 32759
rect 26157 32725 26191 32759
rect 29009 32725 29043 32759
rect 32137 32725 32171 32759
rect 32505 32725 32539 32759
rect 40801 32725 40835 32759
rect 46397 32725 46431 32759
rect 29745 32521 29779 32555
rect 32505 32521 32539 32555
rect 35725 32521 35759 32555
rect 37289 32521 37323 32555
rect 37933 32521 37967 32555
rect 39221 32521 39255 32555
rect 39589 32521 39623 32555
rect 40877 32521 40911 32555
rect 41429 32521 41463 32555
rect 43729 32521 43763 32555
rect 32137 32453 32171 32487
rect 32321 32453 32355 32487
rect 40233 32453 40267 32487
rect 2145 32385 2179 32419
rect 25329 32385 25363 32419
rect 28549 32385 28583 32419
rect 29034 32385 29068 32419
rect 29653 32385 29687 32419
rect 29837 32385 29871 32419
rect 30849 32385 30883 32419
rect 35541 32385 35575 32419
rect 35725 32385 35759 32419
rect 36369 32385 36403 32419
rect 36553 32385 36587 32419
rect 37749 32385 37783 32419
rect 38577 32385 38611 32419
rect 39405 32385 39439 32419
rect 39681 32385 39715 32419
rect 40141 32385 40175 32419
rect 40325 32385 40359 32419
rect 40785 32385 40819 32419
rect 40969 32385 41003 32419
rect 41613 32385 41647 32419
rect 42441 32385 42475 32419
rect 43545 32385 43579 32419
rect 44373 32385 44407 32419
rect 47777 32385 47811 32419
rect 2329 32317 2363 32351
rect 2789 32317 2823 32351
rect 28825 32317 28859 32351
rect 28917 32317 28951 32351
rect 36461 32317 36495 32351
rect 36645 32317 36679 32351
rect 37657 32317 37691 32351
rect 38393 32317 38427 32351
rect 38761 32317 38795 32351
rect 42533 32317 42567 32351
rect 43361 32317 43395 32351
rect 29193 32249 29227 32283
rect 25145 32181 25179 32215
rect 30941 32181 30975 32215
rect 36185 32181 36219 32215
rect 44189 32181 44223 32215
rect 47593 32181 47627 32215
rect 2513 31977 2547 32011
rect 26065 31977 26099 32011
rect 33241 31977 33275 32011
rect 36185 31977 36219 32011
rect 37565 31977 37599 32011
rect 42809 31977 42843 32011
rect 29837 31909 29871 31943
rect 30757 31909 30791 31943
rect 33793 31909 33827 31943
rect 37933 31909 37967 31943
rect 42165 31909 42199 31943
rect 24685 31841 24719 31875
rect 27629 31841 27663 31875
rect 29561 31841 29595 31875
rect 30941 31841 30975 31875
rect 35909 31841 35943 31875
rect 38025 31841 38059 31875
rect 39957 31841 39991 31875
rect 40417 31841 40451 31875
rect 46489 31841 46523 31875
rect 48145 31841 48179 31875
rect 2421 31773 2455 31807
rect 24952 31773 24986 31807
rect 27813 31773 27847 31807
rect 28457 31773 28491 31807
rect 28641 31773 28675 31807
rect 28917 31773 28951 31807
rect 30481 31773 30515 31807
rect 32229 31773 32263 31807
rect 32321 31773 32355 31807
rect 32413 31773 32447 31807
rect 32597 31773 32631 31807
rect 33149 31773 33183 31807
rect 33793 31773 33827 31807
rect 34069 31773 34103 31807
rect 35817 31773 35851 31807
rect 36645 31773 36679 31807
rect 36829 31773 36863 31807
rect 37105 31773 37139 31807
rect 37749 31773 37783 31807
rect 40049 31773 40083 31807
rect 41429 31773 41463 31807
rect 42349 31773 42383 31807
rect 42993 31773 43027 31807
rect 46305 31773 46339 31807
rect 28825 31705 28859 31739
rect 38485 31705 38519 31739
rect 38669 31705 38703 31739
rect 43637 31705 43671 31739
rect 43821 31705 43855 31739
rect 27997 31637 28031 31671
rect 30021 31637 30055 31671
rect 31953 31637 31987 31671
rect 33977 31637 34011 31671
rect 37013 31637 37047 31671
rect 38853 31637 38887 31671
rect 41245 31637 41279 31671
rect 43913 31637 43947 31671
rect 44005 31637 44039 31671
rect 44189 31637 44223 31671
rect 26433 31433 26467 31467
rect 34897 31433 34931 31467
rect 36737 31433 36771 31467
rect 45201 31433 45235 31467
rect 46857 31433 46891 31467
rect 47961 31433 47995 31467
rect 33784 31365 33818 31399
rect 36369 31365 36403 31399
rect 36553 31365 36587 31399
rect 40776 31365 40810 31399
rect 44088 31365 44122 31399
rect 46489 31365 46523 31399
rect 46765 31365 46799 31399
rect 23857 31297 23891 31331
rect 24041 31297 24075 31331
rect 25053 31297 25087 31331
rect 25309 31297 25343 31331
rect 28641 31297 28675 31331
rect 28825 31297 28859 31331
rect 29193 31297 29227 31331
rect 30021 31297 30055 31331
rect 30113 31297 30147 31331
rect 30297 31297 30331 31331
rect 30389 31297 30423 31331
rect 33517 31297 33551 31331
rect 38669 31297 38703 31331
rect 38761 31297 38795 31331
rect 38853 31297 38887 31331
rect 39037 31297 39071 31331
rect 42901 31297 42935 31331
rect 43177 31297 43211 31331
rect 45753 31297 45787 31331
rect 45845 31297 45879 31331
rect 46673 31297 46707 31331
rect 47777 31297 47811 31331
rect 28917 31229 28951 31263
rect 29009 31229 29043 31263
rect 40509 31229 40543 31263
rect 43085 31229 43119 31263
rect 43821 31229 43855 31263
rect 47593 31229 47627 31263
rect 46029 31161 46063 31195
rect 24225 31093 24259 31127
rect 29377 31093 29411 31127
rect 29837 31093 29871 31127
rect 38393 31093 38427 31127
rect 41889 31093 41923 31127
rect 43177 31093 43211 31127
rect 43361 31093 43395 31127
rect 47041 31093 47075 31127
rect 24685 30889 24719 30923
rect 28733 30889 28767 30923
rect 34069 30889 34103 30923
rect 34713 30889 34747 30923
rect 41521 30889 41555 30923
rect 42349 30889 42383 30923
rect 43361 30889 43395 30923
rect 46029 30889 46063 30923
rect 48145 30889 48179 30923
rect 43821 30821 43855 30855
rect 41981 30753 42015 30787
rect 45937 30753 45971 30787
rect 46765 30753 46799 30787
rect 24869 30685 24903 30719
rect 28457 30685 28491 30719
rect 28549 30685 28583 30719
rect 28825 30685 28859 30719
rect 32137 30685 32171 30719
rect 32393 30685 32427 30719
rect 33977 30685 34011 30719
rect 34897 30685 34931 30719
rect 35173 30685 35207 30719
rect 40325 30685 40359 30719
rect 41153 30685 41187 30719
rect 41337 30685 41371 30719
rect 42165 30685 42199 30719
rect 43085 30685 43119 30719
rect 43177 30685 43211 30719
rect 44005 30685 44039 30719
rect 44189 30685 44223 30719
rect 44465 30685 44499 30719
rect 45385 30685 45419 30719
rect 46121 30685 46155 30719
rect 47032 30685 47066 30719
rect 35081 30617 35115 30651
rect 36369 30617 36403 30651
rect 38117 30617 38151 30651
rect 44097 30617 44131 30651
rect 44327 30617 44361 30651
rect 45017 30617 45051 30651
rect 45201 30617 45235 30651
rect 45845 30617 45879 30651
rect 28273 30549 28307 30583
rect 33517 30549 33551 30583
rect 40417 30549 40451 30583
rect 46305 30549 46339 30583
rect 47041 30345 47075 30379
rect 31125 30277 31159 30311
rect 41429 30277 41463 30311
rect 29285 30209 29319 30243
rect 29469 30209 29503 30243
rect 36369 30209 36403 30243
rect 36461 30209 36495 30243
rect 36553 30209 36587 30243
rect 36737 30209 36771 30243
rect 37289 30209 37323 30243
rect 37473 30209 37507 30243
rect 37565 30209 37599 30243
rect 37703 30209 37737 30243
rect 38761 30209 38795 30243
rect 39017 30209 39051 30243
rect 42441 30209 42475 30243
rect 42697 30209 42731 30243
rect 45928 30209 45962 30243
rect 47777 30209 47811 30243
rect 45661 30141 45695 30175
rect 31309 30073 31343 30107
rect 40141 30073 40175 30107
rect 41613 30073 41647 30107
rect 47593 30073 47627 30107
rect 29285 30005 29319 30039
rect 36093 30005 36127 30039
rect 37841 30005 37875 30039
rect 43821 30005 43855 30039
rect 40509 29801 40543 29835
rect 43453 29801 43487 29835
rect 34713 29733 34747 29767
rect 30021 29665 30055 29699
rect 36185 29665 36219 29699
rect 38669 29665 38703 29699
rect 24685 29597 24719 29631
rect 24774 29594 24808 29628
rect 24874 29597 24908 29631
rect 25053 29597 25087 29631
rect 25605 29597 25639 29631
rect 28733 29597 28767 29631
rect 29009 29597 29043 29631
rect 30113 29597 30147 29631
rect 30941 29597 30975 29631
rect 33057 29597 33091 29631
rect 33149 29597 33183 29631
rect 33241 29597 33275 29631
rect 33425 29597 33459 29631
rect 33977 29597 34011 29631
rect 34897 29597 34931 29631
rect 35173 29597 35207 29631
rect 36441 29597 36475 29631
rect 38393 29597 38427 29631
rect 38577 29597 38611 29631
rect 38761 29597 38795 29631
rect 38945 29597 38979 29631
rect 39129 29597 39163 29631
rect 39854 29597 39888 29631
rect 39985 29597 40019 29631
rect 40371 29597 40405 29631
rect 44189 29597 44223 29631
rect 46305 29597 46339 29631
rect 25872 29529 25906 29563
rect 28917 29529 28951 29563
rect 31208 29529 31242 29563
rect 32781 29529 32815 29563
rect 34161 29529 34195 29563
rect 40141 29529 40175 29563
rect 40233 29529 40267 29563
rect 42625 29529 42659 29563
rect 43361 29529 43395 29563
rect 46489 29529 46523 29563
rect 48145 29529 48179 29563
rect 24409 29461 24443 29495
rect 26985 29461 27019 29495
rect 28549 29461 28583 29495
rect 30481 29461 30515 29495
rect 32321 29461 32355 29495
rect 35081 29461 35115 29495
rect 37565 29461 37599 29495
rect 42717 29461 42751 29495
rect 44005 29461 44039 29495
rect 25237 29257 25271 29291
rect 25697 29257 25731 29291
rect 30021 29257 30055 29291
rect 31125 29257 31159 29291
rect 33333 29257 33367 29291
rect 35357 29257 35391 29291
rect 41153 29257 41187 29291
rect 43453 29257 43487 29291
rect 45293 29257 45327 29291
rect 18337 29189 18371 29223
rect 33793 29189 33827 29223
rect 34989 29189 35023 29223
rect 44180 29189 44214 29223
rect 17785 29121 17819 29155
rect 22845 29121 22879 29155
rect 23857 29121 23891 29155
rect 24124 29121 24158 29155
rect 25927 29121 25961 29155
rect 26078 29124 26112 29158
rect 26178 29121 26212 29155
rect 26341 29121 26375 29155
rect 27445 29121 27479 29155
rect 28089 29121 28123 29155
rect 28345 29121 28379 29155
rect 29929 29121 29963 29155
rect 30113 29121 30147 29155
rect 30941 29121 30975 29155
rect 31125 29121 31159 29155
rect 33149 29121 33183 29155
rect 33333 29121 33367 29155
rect 33977 29121 34011 29155
rect 34069 29121 34103 29155
rect 34327 29121 34361 29155
rect 34805 29121 34839 29155
rect 35081 29121 35115 29155
rect 35173 29121 35207 29155
rect 36369 29121 36403 29155
rect 36461 29121 36495 29155
rect 36737 29121 36771 29155
rect 37289 29121 37323 29155
rect 37565 29121 37599 29155
rect 40141 29121 40175 29155
rect 41061 29121 41095 29155
rect 43177 29121 43211 29155
rect 43269 29121 43303 29155
rect 47777 29121 47811 29155
rect 22661 29053 22695 29087
rect 36645 29053 36679 29087
rect 43913 29053 43947 29087
rect 23029 28985 23063 29019
rect 34253 28985 34287 29019
rect 40601 28985 40635 29019
rect 27537 28917 27571 28951
rect 29469 28917 29503 28951
rect 36185 28917 36219 28951
rect 40233 28917 40267 28951
rect 19993 28713 20027 28747
rect 23765 28713 23799 28747
rect 26617 28713 26651 28747
rect 28089 28713 28123 28747
rect 34069 28713 34103 28747
rect 36737 28713 36771 28747
rect 37749 28713 37783 28747
rect 38393 28713 38427 28747
rect 41061 28713 41095 28747
rect 44005 28713 44039 28747
rect 23213 28645 23247 28679
rect 35265 28645 35299 28679
rect 18521 28577 18555 28611
rect 22937 28577 22971 28611
rect 24685 28577 24719 28611
rect 26433 28577 26467 28611
rect 33977 28577 34011 28611
rect 34161 28577 34195 28611
rect 43177 28577 43211 28611
rect 46305 28577 46339 28611
rect 16865 28509 16899 28543
rect 22017 28509 22051 28543
rect 22845 28509 22879 28543
rect 23673 28509 23707 28543
rect 23857 28509 23891 28543
rect 24409 28509 24443 28543
rect 26341 28509 26375 28543
rect 27445 28509 27479 28543
rect 28365 28509 28399 28543
rect 28457 28509 28491 28543
rect 28549 28509 28583 28543
rect 28733 28509 28767 28543
rect 33885 28509 33919 28543
rect 34713 28509 34747 28543
rect 35081 28509 35115 28543
rect 36921 28509 36955 28543
rect 37197 28509 37231 28543
rect 37657 28509 37691 28543
rect 38301 28509 38335 28543
rect 40509 28509 40543 28543
rect 40969 28509 41003 28543
rect 43361 28509 43395 28543
rect 43545 28509 43579 28543
rect 44189 28509 44223 28543
rect 17141 28441 17175 28475
rect 17785 28441 17819 28475
rect 19717 28441 19751 28475
rect 25973 28441 26007 28475
rect 34897 28441 34931 28475
rect 34989 28441 35023 28475
rect 37105 28441 37139 28475
rect 40325 28441 40359 28475
rect 46489 28441 46523 28475
rect 48145 28441 48179 28475
rect 22109 28373 22143 28407
rect 27537 28373 27571 28407
rect 22845 28169 22879 28203
rect 23673 28169 23707 28203
rect 27353 28169 27387 28203
rect 28273 28169 28307 28203
rect 28917 28169 28951 28203
rect 33977 28169 34011 28203
rect 35265 28169 35299 28203
rect 40601 28169 40635 28203
rect 45845 28169 45879 28203
rect 18153 28101 18187 28135
rect 32321 28101 32355 28135
rect 43444 28101 43478 28135
rect 17049 28033 17083 28067
rect 17233 28033 17267 28067
rect 17785 28033 17819 28067
rect 22477 28033 22511 28067
rect 23489 28033 23523 28067
rect 23765 28033 23799 28067
rect 25605 28033 25639 28067
rect 26985 28033 27019 28067
rect 27169 28033 27203 28067
rect 28641 28033 28675 28067
rect 29469 28033 29503 28067
rect 31309 28033 31343 28067
rect 31585 28033 31619 28067
rect 32137 28033 32171 28067
rect 32413 28033 32447 28067
rect 33885 28033 33919 28067
rect 35173 28033 35207 28067
rect 40417 28033 40451 28067
rect 40693 28033 40727 28067
rect 41153 28033 41187 28067
rect 41337 28033 41371 28067
rect 45753 28033 45787 28067
rect 46397 28033 46431 28067
rect 22569 27965 22603 27999
rect 25973 27965 26007 27999
rect 26065 27965 26099 27999
rect 28733 27965 28767 27999
rect 43177 27965 43211 27999
rect 32137 27897 32171 27931
rect 23305 27829 23339 27863
rect 26249 27829 26283 27863
rect 29561 27829 29595 27863
rect 31125 27829 31159 27863
rect 31493 27829 31527 27863
rect 40417 27829 40451 27863
rect 41153 27829 41187 27863
rect 44557 27829 44591 27863
rect 46489 27829 46523 27863
rect 47777 27829 47811 27863
rect 26157 27625 26191 27659
rect 28917 27625 28951 27659
rect 33977 27625 34011 27659
rect 38301 27625 38335 27659
rect 40049 27625 40083 27659
rect 24961 27557 24995 27591
rect 29929 27557 29963 27591
rect 38485 27557 38519 27591
rect 39957 27557 39991 27591
rect 25237 27489 25271 27523
rect 25329 27489 25363 27523
rect 34805 27489 34839 27523
rect 34989 27489 35023 27523
rect 37381 27489 37415 27523
rect 37473 27489 37507 27523
rect 39037 27489 39071 27523
rect 40141 27489 40175 27523
rect 46305 27489 46339 27523
rect 46489 27489 46523 27523
rect 46857 27489 46891 27523
rect 15945 27421 15979 27455
rect 18061 27421 18095 27455
rect 25145 27421 25179 27455
rect 25421 27421 25455 27455
rect 26065 27421 26099 27455
rect 26249 27421 26283 27455
rect 28825 27421 28859 27455
rect 29009 27421 29043 27455
rect 30849 27421 30883 27455
rect 33885 27421 33919 27455
rect 34713 27421 34747 27455
rect 35449 27421 35483 27455
rect 35633 27421 35667 27455
rect 37197 27421 37231 27455
rect 38945 27421 38979 27455
rect 39865 27421 39899 27455
rect 40693 27421 40727 27455
rect 40785 27421 40819 27455
rect 41429 27421 41463 27455
rect 16129 27353 16163 27387
rect 16589 27353 16623 27387
rect 17325 27353 17359 27387
rect 18613 27353 18647 27387
rect 29561 27353 29595 27387
rect 29745 27353 29779 27387
rect 31116 27353 31150 27387
rect 34989 27353 35023 27387
rect 38117 27353 38151 27387
rect 39221 27353 39255 27387
rect 41674 27353 41708 27387
rect 43361 27353 43395 27387
rect 32229 27285 32263 27319
rect 35541 27285 35575 27319
rect 37013 27285 37047 27319
rect 38317 27285 38351 27319
rect 38945 27285 38979 27319
rect 40969 27285 41003 27319
rect 42809 27285 42843 27319
rect 43453 27285 43487 27319
rect 42901 27081 42935 27115
rect 46949 27081 46983 27115
rect 7849 27013 7883 27047
rect 18337 27013 18371 27047
rect 34428 27013 34462 27047
rect 37473 27013 37507 27047
rect 44088 27013 44122 27047
rect 16957 26945 16991 26979
rect 18061 26945 18095 26979
rect 23213 26945 23247 26979
rect 24777 26945 24811 26979
rect 26065 26945 26099 26979
rect 27445 26945 27479 26979
rect 28641 26945 28675 26979
rect 28733 26945 28767 26979
rect 32873 26945 32907 26979
rect 34161 26945 34195 26979
rect 37289 26945 37323 26979
rect 37565 26945 37599 26979
rect 38025 26945 38059 26979
rect 38292 26945 38326 26979
rect 39865 26945 39899 26979
rect 40132 26945 40166 26979
rect 42809 26945 42843 26979
rect 45937 26945 45971 26979
rect 46857 26945 46891 26979
rect 47777 26945 47811 26979
rect 17509 26877 17543 26911
rect 23121 26877 23155 26911
rect 24869 26877 24903 26911
rect 25973 26877 26007 26911
rect 28365 26877 28399 26911
rect 28549 26877 28583 26911
rect 28825 26877 28859 26911
rect 33149 26877 33183 26911
rect 43821 26877 43855 26911
rect 23581 26809 23615 26843
rect 25145 26809 25179 26843
rect 26433 26809 26467 26843
rect 27629 26809 27663 26843
rect 32965 26809 32999 26843
rect 37289 26809 37323 26843
rect 41245 26809 41279 26843
rect 7941 26741 7975 26775
rect 32873 26741 32907 26775
rect 35541 26741 35575 26775
rect 39405 26741 39439 26775
rect 45201 26741 45235 26775
rect 46029 26741 46063 26775
rect 25605 26537 25639 26571
rect 25973 26537 26007 26571
rect 26801 26537 26835 26571
rect 28733 26537 28767 26571
rect 40417 26537 40451 26571
rect 40785 26537 40819 26571
rect 45661 26537 45695 26571
rect 33701 26469 33735 26503
rect 35081 26469 35115 26503
rect 36001 26469 36035 26503
rect 37841 26469 37875 26503
rect 38301 26469 38335 26503
rect 8217 26401 8251 26435
rect 16957 26401 16991 26435
rect 23213 26401 23247 26435
rect 28365 26401 28399 26435
rect 34713 26401 34747 26435
rect 40877 26401 40911 26435
rect 43361 26401 43395 26435
rect 46305 26401 46339 26435
rect 47041 26401 47075 26435
rect 7481 26333 7515 26367
rect 16681 26333 16715 26367
rect 23029 26333 23063 26367
rect 25789 26333 25823 26367
rect 26065 26333 26099 26367
rect 26709 26333 26743 26367
rect 28457 26333 28491 26367
rect 32321 26333 32355 26367
rect 34897 26333 34931 26367
rect 36461 26333 36495 26367
rect 38577 26333 38611 26367
rect 40601 26333 40635 26367
rect 45017 26333 45051 26367
rect 45293 26333 45327 26367
rect 45385 26333 45419 26367
rect 46121 26333 46155 26367
rect 32588 26265 32622 26299
rect 35817 26265 35851 26299
rect 36728 26265 36762 26299
rect 38301 26265 38335 26299
rect 41613 26265 41647 26299
rect 45502 26265 45536 26299
rect 38485 26197 38519 26231
rect 26249 25993 26283 26027
rect 27077 25993 27111 26027
rect 28641 25993 28675 26027
rect 29929 25993 29963 26027
rect 33793 25993 33827 26027
rect 40325 25993 40359 26027
rect 29561 25925 29595 25959
rect 29761 25925 29795 25959
rect 32689 25925 32723 25959
rect 33425 25925 33459 25959
rect 33625 25925 33659 25959
rect 45845 25925 45879 25959
rect 8033 25857 8067 25891
rect 9229 25857 9263 25891
rect 22201 25857 22235 25891
rect 25136 25857 25170 25891
rect 26985 25857 27019 25891
rect 27997 25857 28031 25891
rect 28181 25857 28215 25891
rect 28825 25857 28859 25891
rect 30573 25857 30607 25891
rect 30757 25857 30791 25891
rect 31125 25857 31159 25891
rect 32873 25857 32907 25891
rect 32965 25857 32999 25891
rect 36461 25857 36495 25891
rect 39037 25857 39071 25891
rect 43637 25857 43671 25891
rect 45477 25857 45511 25891
rect 45661 25857 45695 25891
rect 46305 25857 46339 25891
rect 46489 25857 46523 25891
rect 47593 25857 47627 25891
rect 8585 25789 8619 25823
rect 9505 25789 9539 25823
rect 22293 25789 22327 25823
rect 24869 25789 24903 25823
rect 29101 25789 29135 25823
rect 30849 25789 30883 25823
rect 30941 25789 30975 25823
rect 44557 25789 44591 25823
rect 32689 25721 32723 25755
rect 44005 25721 44039 25755
rect 44833 25721 44867 25755
rect 46305 25721 46339 25755
rect 22477 25653 22511 25687
rect 28089 25653 28123 25687
rect 29009 25653 29043 25687
rect 29745 25653 29779 25687
rect 31309 25653 31343 25687
rect 33609 25653 33643 25687
rect 36553 25653 36587 25687
rect 44097 25653 44131 25687
rect 45017 25653 45051 25687
rect 47685 25653 47719 25687
rect 25513 25449 25547 25483
rect 32137 25449 32171 25483
rect 40417 25449 40451 25483
rect 44373 25449 44407 25483
rect 25421 25381 25455 25415
rect 26065 25381 26099 25415
rect 29653 25381 29687 25415
rect 35817 25381 35851 25415
rect 46489 25313 46523 25347
rect 46765 25313 46799 25347
rect 2145 25245 2179 25279
rect 2605 25245 2639 25279
rect 7849 25245 7883 25279
rect 8125 25245 8159 25279
rect 21833 25245 21867 25279
rect 22017 25245 22051 25279
rect 22477 25245 22511 25279
rect 22661 25245 22695 25279
rect 23305 25245 23339 25279
rect 23489 25245 23523 25279
rect 25145 25245 25179 25279
rect 25329 25245 25363 25279
rect 25513 25245 25547 25279
rect 26065 25245 26099 25279
rect 26249 25245 26283 25279
rect 27905 25245 27939 25279
rect 28733 25245 28767 25279
rect 28917 25245 28951 25279
rect 29009 25245 29043 25279
rect 29561 25245 29595 25279
rect 30757 25245 30791 25279
rect 35817 25245 35851 25279
rect 36001 25245 36035 25279
rect 40969 25245 41003 25279
rect 44097 25245 44131 25279
rect 44189 25245 44223 25279
rect 44465 25245 44499 25279
rect 45201 25245 45235 25279
rect 45385 25245 45419 25279
rect 45477 25245 45511 25279
rect 46305 25245 46339 25279
rect 31024 25177 31058 25211
rect 40325 25177 40359 25211
rect 2697 25109 2731 25143
rect 22017 25109 22051 25143
rect 22845 25109 22879 25143
rect 23397 25109 23431 25143
rect 27997 25109 28031 25143
rect 28549 25109 28583 25143
rect 41061 25109 41095 25143
rect 43913 25109 43947 25143
rect 45017 25109 45051 25143
rect 28181 24905 28215 24939
rect 2329 24837 2363 24871
rect 2145 24769 2179 24803
rect 7849 24769 7883 24803
rect 24777 24769 24811 24803
rect 27813 24769 27847 24803
rect 28641 24769 28675 24803
rect 28825 24769 28859 24803
rect 31033 24769 31067 24803
rect 35817 24769 35851 24803
rect 36461 24769 36495 24803
rect 38025 24769 38059 24803
rect 38292 24769 38326 24803
rect 39865 24769 39899 24803
rect 40049 24769 40083 24803
rect 44005 24769 44039 24803
rect 44189 24769 44223 24803
rect 44281 24769 44315 24803
rect 44557 24769 44591 24803
rect 45385 24769 45419 24803
rect 45477 24769 45511 24803
rect 45661 24769 45695 24803
rect 45753 24769 45787 24803
rect 46305 24769 46339 24803
rect 47777 24769 47811 24803
rect 2789 24701 2823 24735
rect 8033 24701 8067 24735
rect 22017 24701 22051 24735
rect 22201 24701 22235 24735
rect 22477 24701 22511 24735
rect 27905 24701 27939 24735
rect 28733 24701 28767 24735
rect 33333 24701 33367 24735
rect 33609 24701 33643 24735
rect 35633 24701 35667 24735
rect 36737 24701 36771 24735
rect 44373 24701 44407 24735
rect 36645 24633 36679 24667
rect 24869 24565 24903 24599
rect 31125 24565 31159 24599
rect 36001 24565 36035 24599
rect 36553 24565 36587 24599
rect 39405 24565 39439 24599
rect 39865 24565 39899 24599
rect 44741 24565 44775 24599
rect 45201 24565 45235 24599
rect 46397 24565 46431 24599
rect 22109 24361 22143 24395
rect 23305 24361 23339 24395
rect 38025 24361 38059 24395
rect 39037 24361 39071 24395
rect 39865 24361 39899 24395
rect 30481 24225 30515 24259
rect 35541 24225 35575 24259
rect 38209 24225 38243 24259
rect 41429 24225 41463 24259
rect 43085 24225 43119 24259
rect 46305 24225 46339 24259
rect 48145 24225 48179 24259
rect 2329 24157 2363 24191
rect 22017 24157 22051 24191
rect 22937 24157 22971 24191
rect 23397 24157 23431 24191
rect 24409 24157 24443 24191
rect 27629 24157 27663 24191
rect 30389 24157 30423 24191
rect 31493 24157 31527 24191
rect 31585 24157 31619 24191
rect 31769 24157 31803 24191
rect 31861 24157 31895 24191
rect 32965 24157 32999 24191
rect 33149 24157 33183 24191
rect 33241 24157 33275 24191
rect 33885 24157 33919 24191
rect 33977 24157 34011 24191
rect 34897 24157 34931 24191
rect 35081 24157 35115 24191
rect 35808 24157 35842 24191
rect 37933 24157 37967 24191
rect 38761 24157 38795 24191
rect 38853 24157 38887 24191
rect 39865 24157 39899 24191
rect 40049 24157 40083 24191
rect 41245 24157 41279 24191
rect 43821 24157 43855 24191
rect 44005 24157 44039 24191
rect 45201 24157 45235 24191
rect 45477 24157 45511 24191
rect 23029 24089 23063 24123
rect 24654 24089 24688 24123
rect 27813 24089 27847 24123
rect 33701 24089 33735 24123
rect 38209 24089 38243 24123
rect 45385 24089 45419 24123
rect 46489 24089 46523 24123
rect 23121 24021 23155 24055
rect 23397 24021 23431 24055
rect 25789 24021 25823 24055
rect 27997 24021 28031 24055
rect 31309 24021 31343 24055
rect 32781 24021 32815 24055
rect 33799 24021 33833 24055
rect 34989 24021 35023 24055
rect 36921 24021 36955 24055
rect 43913 24021 43947 24055
rect 45017 24021 45051 24055
rect 24041 23817 24075 23851
rect 33885 23817 33919 23851
rect 36553 23817 36587 23851
rect 38685 23817 38719 23851
rect 38853 23817 38887 23851
rect 39589 23817 39623 23851
rect 43177 23817 43211 23851
rect 46949 23817 46983 23851
rect 27721 23749 27755 23783
rect 28641 23749 28675 23783
rect 32772 23749 32806 23783
rect 36185 23749 36219 23783
rect 36401 23749 36435 23783
rect 38485 23749 38519 23783
rect 2053 23681 2087 23715
rect 24409 23681 24443 23715
rect 24777 23681 24811 23715
rect 25421 23681 25455 23715
rect 25514 23681 25548 23715
rect 25697 23681 25731 23715
rect 25786 23681 25820 23715
rect 25925 23681 25959 23715
rect 26985 23681 27019 23715
rect 27169 23683 27203 23717
rect 27537 23681 27571 23715
rect 30849 23681 30883 23715
rect 31033 23681 31067 23715
rect 31125 23681 31159 23715
rect 31401 23681 31435 23715
rect 32505 23681 32539 23715
rect 34345 23681 34379 23715
rect 34612 23681 34646 23715
rect 39313 23681 39347 23715
rect 40509 23681 40543 23715
rect 40765 23681 40799 23715
rect 43085 23681 43119 23715
rect 43269 23681 43303 23715
rect 43913 23681 43947 23715
rect 45891 23681 45925 23715
rect 46029 23681 46063 23715
rect 46121 23681 46155 23715
rect 46305 23681 46339 23715
rect 46857 23681 46891 23715
rect 47777 23681 47811 23715
rect 2237 23613 2271 23647
rect 2789 23613 2823 23647
rect 23949 23613 23983 23647
rect 24317 23613 24351 23647
rect 24685 23613 24719 23647
rect 27255 23613 27289 23647
rect 27353 23613 27387 23647
rect 31217 23613 31251 23647
rect 39589 23613 39623 23647
rect 43821 23613 43855 23647
rect 26065 23545 26099 23579
rect 39405 23545 39439 23579
rect 44281 23545 44315 23579
rect 29929 23477 29963 23511
rect 31585 23477 31619 23511
rect 35725 23477 35759 23511
rect 36369 23477 36403 23511
rect 38669 23477 38703 23511
rect 41889 23477 41923 23511
rect 45661 23477 45695 23511
rect 2421 23273 2455 23307
rect 24409 23273 24443 23307
rect 27813 23273 27847 23307
rect 32505 23273 32539 23307
rect 35081 23273 35115 23307
rect 35449 23273 35483 23307
rect 41337 23273 41371 23307
rect 45109 23273 45143 23307
rect 48053 23273 48087 23307
rect 24869 23205 24903 23239
rect 29009 23205 29043 23239
rect 30481 23205 30515 23239
rect 2329 23069 2363 23103
rect 24593 23069 24627 23103
rect 24685 23069 24719 23103
rect 24961 23069 24995 23103
rect 27261 23069 27295 23103
rect 27445 23069 27479 23103
rect 27629 23069 27663 23103
rect 28365 23069 28399 23103
rect 28513 23069 28547 23103
rect 28733 23069 28767 23103
rect 28830 23069 28864 23103
rect 30757 23069 30791 23103
rect 31217 23069 31251 23103
rect 35265 23069 35299 23103
rect 35541 23069 35575 23103
rect 36277 23069 36311 23103
rect 37749 23069 37783 23103
rect 39865 23069 39899 23103
rect 40601 23069 40635 23103
rect 40785 23069 40819 23103
rect 40877 23069 40911 23103
rect 40969 23069 41003 23103
rect 41153 23069 41187 23103
rect 45017 23069 45051 23103
rect 45201 23069 45235 23103
rect 46673 23069 46707 23103
rect 46940 23069 46974 23103
rect 27537 23001 27571 23035
rect 28641 23001 28675 23035
rect 30481 23001 30515 23035
rect 30665 22933 30699 22967
rect 36369 22933 36403 22967
rect 37841 22933 37875 22967
rect 39957 22933 39991 22967
rect 30941 22729 30975 22763
rect 34437 22729 34471 22763
rect 38025 22729 38059 22763
rect 39865 22729 39899 22763
rect 41061 22729 41095 22763
rect 24409 22661 24443 22695
rect 32505 22661 32539 22695
rect 33302 22661 33336 22695
rect 35909 22661 35943 22695
rect 36093 22661 36127 22695
rect 39497 22661 39531 22695
rect 45477 22661 45511 22695
rect 24593 22593 24627 22627
rect 24685 22593 24719 22627
rect 29561 22593 29595 22627
rect 29828 22593 29862 22627
rect 31585 22593 31619 22627
rect 32413 22593 32447 22627
rect 32597 22593 32631 22627
rect 36185 22593 36219 22627
rect 37289 22593 37323 22627
rect 37933 22593 37967 22627
rect 38669 22593 38703 22627
rect 39313 22593 39347 22627
rect 39589 22593 39623 22627
rect 39681 22593 39715 22627
rect 40325 22593 40359 22627
rect 40509 22593 40543 22627
rect 40693 22593 40727 22627
rect 40877 22593 40911 22627
rect 42441 22593 42475 22627
rect 42697 22593 42731 22627
rect 45293 22593 45327 22627
rect 47593 22593 47627 22627
rect 33057 22525 33091 22559
rect 40601 22525 40635 22559
rect 37381 22457 37415 22491
rect 24409 22389 24443 22423
rect 31401 22389 31435 22423
rect 35909 22389 35943 22423
rect 38761 22389 38795 22423
rect 43821 22389 43855 22423
rect 45661 22389 45695 22423
rect 47041 22389 47075 22423
rect 47685 22389 47719 22423
rect 25789 22185 25823 22219
rect 26433 22185 26467 22219
rect 30021 22185 30055 22219
rect 30389 22185 30423 22219
rect 40601 22185 40635 22219
rect 42441 22185 42475 22219
rect 27353 22049 27387 22083
rect 31033 22049 31067 22083
rect 31309 22049 31343 22083
rect 32597 22049 32631 22083
rect 35817 22049 35851 22083
rect 45293 22049 45327 22083
rect 46305 22049 46339 22083
rect 48145 22049 48179 22083
rect 2329 21981 2363 22015
rect 24409 21981 24443 22015
rect 27077 21981 27111 22015
rect 27169 21981 27203 22015
rect 30205 21981 30239 22015
rect 30481 21981 30515 22015
rect 32321 21981 32355 22015
rect 38945 21981 38979 22015
rect 39957 21981 39991 22015
rect 40050 21981 40084 22015
rect 40422 21981 40456 22015
rect 41705 21981 41739 22015
rect 41889 21981 41923 22015
rect 41981 21981 42015 22015
rect 42073 21981 42107 22015
rect 42257 21981 42291 22015
rect 42901 21981 42935 22015
rect 43085 21981 43119 22015
rect 45201 21981 45235 22015
rect 45385 21981 45419 22015
rect 45477 21981 45511 22015
rect 24676 21913 24710 21947
rect 26249 21913 26283 21947
rect 36062 21913 36096 21947
rect 39129 21913 39163 21947
rect 40233 21913 40267 21947
rect 40325 21913 40359 21947
rect 46489 21913 46523 21947
rect 26449 21845 26483 21879
rect 26617 21845 26651 21879
rect 27353 21845 27387 21879
rect 37197 21845 37231 21879
rect 39313 21845 39347 21879
rect 42993 21845 43027 21879
rect 45017 21845 45051 21879
rect 25145 21641 25179 21675
rect 30405 21641 30439 21675
rect 35909 21641 35943 21675
rect 40233 21641 40267 21675
rect 41889 21641 41923 21675
rect 42993 21641 43027 21675
rect 45017 21641 45051 21675
rect 30205 21573 30239 21607
rect 31033 21573 31067 21607
rect 2053 21505 2087 21539
rect 24317 21505 24351 21539
rect 25053 21505 25087 21539
rect 25237 21505 25271 21539
rect 27169 21505 27203 21539
rect 27905 21505 27939 21539
rect 27997 21505 28031 21539
rect 28641 21505 28675 21539
rect 28825 21505 28859 21539
rect 31217 21505 31251 21539
rect 31309 21505 31343 21539
rect 34437 21505 34471 21539
rect 36093 21505 36127 21539
rect 36277 21505 36311 21539
rect 38301 21505 38335 21539
rect 38485 21505 38519 21539
rect 38669 21505 38703 21539
rect 38853 21505 38887 21539
rect 39497 21505 39531 21539
rect 39681 21505 39715 21539
rect 39865 21505 39899 21539
rect 40049 21505 40083 21539
rect 41705 21505 41739 21539
rect 41889 21505 41923 21539
rect 42809 21505 42843 21539
rect 43085 21505 43119 21539
rect 44189 21505 44223 21539
rect 45385 21505 45419 21539
rect 46213 21505 46247 21539
rect 47777 21505 47811 21539
rect 2237 21437 2271 21471
rect 2789 21437 2823 21471
rect 24593 21437 24627 21471
rect 26985 21437 27019 21471
rect 36369 21437 36403 21471
rect 38577 21437 38611 21471
rect 39037 21437 39071 21471
rect 39773 21437 39807 21471
rect 42625 21437 42659 21471
rect 44281 21437 44315 21471
rect 44557 21437 44591 21471
rect 45477 21437 45511 21471
rect 46489 21437 46523 21471
rect 47685 21437 47719 21471
rect 24501 21369 24535 21403
rect 30573 21369 30607 21403
rect 34529 21369 34563 21403
rect 48145 21369 48179 21403
rect 24133 21301 24167 21335
rect 27353 21301 27387 21335
rect 28181 21301 28215 21335
rect 28641 21301 28675 21335
rect 30389 21301 30423 21335
rect 31033 21301 31067 21335
rect 45661 21301 45695 21335
rect 2421 21097 2455 21131
rect 25789 21097 25823 21131
rect 26985 21097 27019 21131
rect 29009 21097 29043 21131
rect 31309 21097 31343 21131
rect 38117 21097 38151 21131
rect 40417 21097 40451 21131
rect 42993 21097 43027 21131
rect 45109 21097 45143 21131
rect 48145 21097 48179 21131
rect 33701 21029 33735 21063
rect 39037 21029 39071 21063
rect 43177 21029 43211 21063
rect 27169 20961 27203 20995
rect 29929 20961 29963 20995
rect 46765 20961 46799 20995
rect 2329 20893 2363 20927
rect 3157 20893 3191 20927
rect 24409 20893 24443 20927
rect 26249 20893 26283 20927
rect 26433 20893 26467 20927
rect 26893 20893 26927 20927
rect 27629 20893 27663 20927
rect 31769 20893 31803 20927
rect 31953 20893 31987 20927
rect 33885 20893 33919 20927
rect 33977 20893 34011 20927
rect 34897 20893 34931 20927
rect 35173 20893 35207 20927
rect 35633 20893 35667 20927
rect 37473 20893 37507 20927
rect 37621 20893 37655 20927
rect 37938 20893 37972 20927
rect 39037 20893 39071 20927
rect 39313 20893 39347 20927
rect 39865 20893 39899 20927
rect 40233 20893 40267 20927
rect 45017 20893 45051 20927
rect 45201 20893 45235 20927
rect 45891 20893 45925 20927
rect 46029 20893 46063 20927
rect 46121 20893 46155 20927
rect 46305 20893 46339 20927
rect 24654 20825 24688 20859
rect 27896 20825 27930 20859
rect 30196 20825 30230 20859
rect 31861 20825 31895 20859
rect 33701 20825 33735 20859
rect 34713 20825 34747 20859
rect 37749 20825 37783 20859
rect 37841 20825 37875 20859
rect 40049 20825 40083 20859
rect 40141 20825 40175 20859
rect 42809 20825 42843 20859
rect 45661 20825 45695 20859
rect 47010 20825 47044 20859
rect 26341 20757 26375 20791
rect 27169 20757 27203 20791
rect 35081 20757 35115 20791
rect 35725 20757 35759 20791
rect 39221 20757 39255 20791
rect 43009 20757 43043 20791
rect 28457 20553 28491 20587
rect 31309 20553 31343 20587
rect 35725 20553 35759 20587
rect 37289 20553 37323 20587
rect 44649 20553 44683 20587
rect 27353 20485 27387 20519
rect 27569 20485 27603 20519
rect 33057 20485 33091 20519
rect 2145 20417 2179 20451
rect 26065 20417 26099 20451
rect 26341 20417 26375 20451
rect 28181 20417 28215 20451
rect 29929 20417 29963 20451
rect 30196 20417 30230 20451
rect 33241 20417 33275 20451
rect 33333 20417 33367 20451
rect 33793 20417 33827 20451
rect 34049 20417 34083 20451
rect 35633 20417 35667 20451
rect 37565 20417 37599 20451
rect 37657 20417 37691 20451
rect 37749 20417 37783 20451
rect 37933 20417 37967 20451
rect 39129 20417 39163 20451
rect 39405 20417 39439 20451
rect 44833 20417 44867 20451
rect 45109 20417 45143 20451
rect 47593 20417 47627 20451
rect 2329 20349 2363 20383
rect 2789 20349 2823 20383
rect 28457 20349 28491 20383
rect 45017 20349 45051 20383
rect 26249 20281 26283 20315
rect 27721 20281 27755 20315
rect 25881 20213 25915 20247
rect 27537 20213 27571 20247
rect 28273 20213 28307 20247
rect 33057 20213 33091 20247
rect 35173 20213 35207 20247
rect 38945 20213 38979 20247
rect 39313 20213 39347 20247
rect 47685 20213 47719 20247
rect 2605 20009 2639 20043
rect 26249 20009 26283 20043
rect 28089 20009 28123 20043
rect 30205 20009 30239 20043
rect 33793 20009 33827 20043
rect 34897 20009 34931 20043
rect 35081 20009 35115 20043
rect 37473 20009 37507 20043
rect 41613 20009 41647 20043
rect 45569 20009 45603 20043
rect 30297 19941 30331 19975
rect 33701 19941 33735 19975
rect 38209 19941 38243 19975
rect 24869 19873 24903 19907
rect 31769 19873 31803 19907
rect 36093 19873 36127 19907
rect 42073 19873 42107 19907
rect 46489 19873 46523 19907
rect 48145 19873 48179 19907
rect 2513 19805 2547 19839
rect 26709 19805 26743 19839
rect 30205 19805 30239 19839
rect 30481 19805 30515 19839
rect 33609 19805 33643 19839
rect 36360 19805 36394 19839
rect 38025 19805 38059 19839
rect 38761 19805 38795 19839
rect 38945 19805 38979 19839
rect 40233 19805 40267 19839
rect 44281 19805 44315 19839
rect 45477 19805 45511 19839
rect 46305 19805 46339 19839
rect 25136 19737 25170 19771
rect 26976 19737 27010 19771
rect 32036 19737 32070 19771
rect 33885 19737 33919 19771
rect 34713 19737 34747 19771
rect 40478 19737 40512 19771
rect 42340 19737 42374 19771
rect 33149 19669 33183 19703
rect 34913 19669 34947 19703
rect 38853 19669 38887 19703
rect 43453 19669 43487 19703
rect 44373 19669 44407 19703
rect 27169 19465 27203 19499
rect 32413 19465 32447 19499
rect 34437 19465 34471 19499
rect 39221 19465 39255 19499
rect 44557 19465 44591 19499
rect 47041 19465 47075 19499
rect 33324 19397 33358 19431
rect 41705 19397 41739 19431
rect 45906 19397 45940 19431
rect 27077 19329 27111 19363
rect 27261 19329 27295 19363
rect 32321 19329 32355 19363
rect 32505 19329 32539 19363
rect 33057 19329 33091 19363
rect 37289 19329 37323 19363
rect 37556 19329 37590 19363
rect 39129 19329 39163 19363
rect 40463 19329 40497 19363
rect 40598 19329 40632 19363
rect 40693 19329 40727 19363
rect 40877 19329 40911 19363
rect 42441 19329 42475 19363
rect 42625 19329 42659 19363
rect 43269 19329 43303 19363
rect 43545 19329 43579 19363
rect 44787 19329 44821 19363
rect 44922 19329 44956 19363
rect 45022 19329 45056 19363
rect 45201 19329 45235 19363
rect 45661 19329 45695 19363
rect 40233 19261 40267 19295
rect 47777 19261 47811 19295
rect 38669 19193 38703 19227
rect 41889 19193 41923 19227
rect 42441 19125 42475 19159
rect 38669 18921 38703 18955
rect 40509 18921 40543 18955
rect 42073 18921 42107 18955
rect 42257 18921 42291 18955
rect 43545 18921 43579 18955
rect 45247 18921 45281 18955
rect 38761 18853 38795 18887
rect 42165 18785 42199 18819
rect 43637 18785 43671 18819
rect 45017 18785 45051 18819
rect 48145 18785 48179 18819
rect 2329 18717 2363 18751
rect 2789 18717 2823 18751
rect 38761 18717 38795 18751
rect 40417 18717 40451 18751
rect 40601 18717 40635 18751
rect 41981 18717 42015 18751
rect 43361 18717 43395 18751
rect 44281 18717 44315 18751
rect 46305 18717 46339 18751
rect 38393 18649 38427 18683
rect 41797 18649 41831 18683
rect 44097 18649 44131 18683
rect 46489 18649 46523 18683
rect 2881 18581 2915 18615
rect 38485 18581 38519 18615
rect 43177 18581 43211 18615
rect 44465 18581 44499 18615
rect 44373 18377 44407 18411
rect 45017 18377 45051 18411
rect 46949 18377 46983 18411
rect 2329 18309 2363 18343
rect 42533 18309 42567 18343
rect 42717 18309 42751 18343
rect 43177 18309 43211 18343
rect 2145 18241 2179 18275
rect 43545 18241 43579 18275
rect 44741 18241 44775 18275
rect 44833 18241 44867 18275
rect 45661 18241 45695 18275
rect 46857 18241 46891 18275
rect 47777 18241 47811 18275
rect 2789 18173 2823 18207
rect 13001 18173 13035 18207
rect 13461 18173 13495 18207
rect 13645 18173 13679 18207
rect 15117 18173 15151 18207
rect 43637 18173 43671 18207
rect 45569 18173 45603 18207
rect 46029 18105 46063 18139
rect 43821 18037 43855 18071
rect 13185 17833 13219 17867
rect 38209 17765 38243 17799
rect 39221 17765 39255 17799
rect 43085 17765 43119 17799
rect 37933 17697 37967 17731
rect 38761 17697 38795 17731
rect 41061 17697 41095 17731
rect 42625 17697 42659 17731
rect 44005 17697 44039 17731
rect 2329 17629 2363 17663
rect 13093 17629 13127 17663
rect 37841 17629 37875 17663
rect 38853 17629 38887 17663
rect 40417 17629 40451 17663
rect 40601 17629 40635 17663
rect 41245 17629 41279 17663
rect 42717 17629 42751 17663
rect 43729 17629 43763 17663
rect 43821 17629 43855 17663
rect 43913 17629 43947 17663
rect 41429 17561 41463 17595
rect 40509 17493 40543 17527
rect 43545 17493 43579 17527
rect 40509 17289 40543 17323
rect 44189 17289 44223 17323
rect 2145 17153 2179 17187
rect 40141 17153 40175 17187
rect 40969 17153 41003 17187
rect 41153 17153 41187 17187
rect 42625 17153 42659 17187
rect 44097 17153 44131 17187
rect 44281 17153 44315 17187
rect 46857 17153 46891 17187
rect 2329 17085 2363 17119
rect 2789 17085 2823 17119
rect 40049 17085 40083 17119
rect 41061 17085 41095 17119
rect 42717 17085 42751 17119
rect 42993 17085 43027 17119
rect 46949 16949 46983 16983
rect 47777 16949 47811 16983
rect 2513 16745 2547 16779
rect 39865 16745 39899 16779
rect 46305 16609 46339 16643
rect 48145 16609 48179 16643
rect 2421 16551 2455 16585
rect 40049 16541 40083 16575
rect 40325 16541 40359 16575
rect 46489 16473 46523 16507
rect 40233 16405 40267 16439
rect 2329 15453 2363 15487
rect 47685 15453 47719 15487
rect 2145 14977 2179 15011
rect 47593 14977 47627 15011
rect 2329 14909 2363 14943
rect 2789 14909 2823 14943
rect 47685 14773 47719 14807
rect 2605 14569 2639 14603
rect 46305 14433 46339 14467
rect 46489 14433 46523 14467
rect 48145 14433 48179 14467
rect 1869 14365 1903 14399
rect 2513 14365 2547 14399
rect 3985 14365 4019 14399
rect 1961 14229 1995 14263
rect 2329 13957 2363 13991
rect 2145 13889 2179 13923
rect 2789 13821 2823 13855
rect 47777 13685 47811 13719
rect 46305 13345 46339 13379
rect 48145 13345 48179 13379
rect 46489 13209 46523 13243
rect 47685 12937 47719 12971
rect 46213 12801 46247 12835
rect 47593 12801 47627 12835
rect 46305 12597 46339 12631
rect 47041 12597 47075 12631
rect 46305 12257 46339 12291
rect 46489 12257 46523 12291
rect 48145 12257 48179 12291
rect 2329 12189 2363 12223
rect 2053 11713 2087 11747
rect 46765 11713 46799 11747
rect 2237 11645 2271 11679
rect 2789 11645 2823 11679
rect 46857 11509 46891 11543
rect 47777 11509 47811 11543
rect 2421 11305 2455 11339
rect 46305 11169 46339 11203
rect 46489 11169 46523 11203
rect 46857 11169 46891 11203
rect 2329 11101 2363 11135
rect 3157 11101 3191 11135
rect 2145 10625 2179 10659
rect 2329 10557 2363 10591
rect 3709 10557 3743 10591
rect 2237 10217 2271 10251
rect 2145 10013 2179 10047
rect 2973 10013 3007 10047
rect 3801 10013 3835 10047
rect 19717 10013 19751 10047
rect 26433 10013 26467 10047
rect 20085 9945 20119 9979
rect 3893 9877 3927 9911
rect 26525 9877 26559 9911
rect 2973 9605 3007 9639
rect 2145 9537 2179 9571
rect 2789 9537 2823 9571
rect 3249 9469 3283 9503
rect 2237 9333 2271 9367
rect 2329 8925 2363 8959
rect 48053 8585 48087 8619
rect 2329 8517 2363 8551
rect 2145 8449 2179 8483
rect 47961 8449 47995 8483
rect 2881 8381 2915 8415
rect 2329 7837 2363 7871
rect 2789 7837 2823 7871
rect 2881 7701 2915 7735
rect 2329 7429 2363 7463
rect 2145 7361 2179 7395
rect 47593 7361 47627 7395
rect 2789 7293 2823 7327
rect 1685 7157 1719 7191
rect 47685 7157 47719 7191
rect 46489 6817 46523 6851
rect 48145 6817 48179 6851
rect 2421 6749 2455 6783
rect 46305 6749 46339 6783
rect 2513 6613 2547 6647
rect 2329 6341 2363 6375
rect 2145 6273 2179 6307
rect 46213 6273 46247 6307
rect 46857 6273 46891 6307
rect 47777 6273 47811 6307
rect 2789 6205 2823 6239
rect 46305 6069 46339 6103
rect 46949 6069 46983 6103
rect 1961 5661 1995 5695
rect 2605 5661 2639 5695
rect 3801 5661 3835 5695
rect 45661 5661 45695 5695
rect 46305 5661 46339 5695
rect 45753 5593 45787 5627
rect 46489 5593 46523 5627
rect 48145 5593 48179 5627
rect 3893 5525 3927 5559
rect 2605 5253 2639 5287
rect 45385 5253 45419 5287
rect 2421 5185 2455 5219
rect 2881 5117 2915 5151
rect 44741 5117 44775 5151
rect 45201 5117 45235 5151
rect 46857 5117 46891 5151
rect 1961 4981 1995 5015
rect 47777 4981 47811 5015
rect 44465 4777 44499 4811
rect 46305 4641 46339 4675
rect 46489 4641 46523 4675
rect 48145 4641 48179 4675
rect 1685 4573 1719 4607
rect 2329 4573 2363 4607
rect 2973 4573 3007 4607
rect 4445 4573 4479 4607
rect 4905 4573 4939 4607
rect 6377 4573 6411 4607
rect 8033 4573 8067 4607
rect 8953 4573 8987 4607
rect 19257 4573 19291 4607
rect 19901 4573 19935 4607
rect 42349 4573 42383 4607
rect 45293 4573 45327 4607
rect 1777 4505 1811 4539
rect 2421 4437 2455 4471
rect 3065 4437 3099 4471
rect 4997 4437 5031 4471
rect 9045 4437 9079 4471
rect 19349 4437 19383 4471
rect 19993 4437 20027 4471
rect 45385 4437 45419 4471
rect 45385 4165 45419 4199
rect 1501 4097 1535 4131
rect 2145 4097 2179 4131
rect 4537 4097 4571 4131
rect 6377 4097 6411 4131
rect 7113 4097 7147 4131
rect 7757 4097 7791 4131
rect 22109 4097 22143 4131
rect 25421 4097 25455 4131
rect 38669 4097 38703 4131
rect 40049 4097 40083 4131
rect 40785 4097 40819 4131
rect 41705 4097 41739 4131
rect 43545 4097 43579 4131
rect 2329 4029 2363 4063
rect 3157 4029 3191 4063
rect 7941 4029 7975 4063
rect 8677 4029 8711 4063
rect 12357 4029 12391 4063
rect 12541 4029 12575 4063
rect 12909 4029 12943 4063
rect 18245 4029 18279 4063
rect 18705 4029 18739 4063
rect 18889 4029 18923 4063
rect 19441 4029 19475 4063
rect 45201 4029 45235 4063
rect 47041 4029 47075 4063
rect 39497 3961 39531 3995
rect 47777 3961 47811 3995
rect 1593 3893 1627 3927
rect 4629 3893 4663 3927
rect 5825 3893 5859 3927
rect 6469 3893 6503 3927
rect 7205 3893 7239 3927
rect 10701 3893 10735 3927
rect 17417 3893 17451 3927
rect 22201 3893 22235 3927
rect 25513 3893 25547 3927
rect 38761 3893 38795 3927
rect 40141 3893 40175 3927
rect 40877 3893 40911 3927
rect 41797 3893 41831 3927
rect 42625 3893 42659 3927
rect 43637 3893 43671 3927
rect 44373 3893 44407 3927
rect 12817 3689 12851 3723
rect 1593 3553 1627 3587
rect 1869 3553 1903 3587
rect 3985 3553 4019 3587
rect 4261 3553 4295 3587
rect 6101 3553 6135 3587
rect 6285 3553 6319 3587
rect 6561 3553 6595 3587
rect 10425 3553 10459 3587
rect 10977 3553 11011 3587
rect 25513 3553 25547 3587
rect 26709 3553 26743 3587
rect 40049 3553 40083 3587
rect 40601 3553 40635 3587
rect 42165 3553 42199 3587
rect 42349 3553 42383 3587
rect 42625 3553 42659 3587
rect 46305 3553 46339 3587
rect 47777 3553 47811 3587
rect 1409 3485 1443 3519
rect 3801 3485 3835 3519
rect 8953 3485 8987 3519
rect 9781 3485 9815 3519
rect 12725 3485 12759 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 17233 3485 17267 3519
rect 17877 3485 17911 3519
rect 18705 3485 18739 3519
rect 19533 3485 19567 3519
rect 22201 3485 22235 3519
rect 25329 3485 25363 3519
rect 27813 3485 27847 3519
rect 28273 3485 28307 3519
rect 31769 3485 31803 3519
rect 32229 3485 32263 3519
rect 39313 3485 39347 3519
rect 39865 3485 39899 3519
rect 45017 3485 45051 3519
rect 45845 3485 45879 3519
rect 10609 3417 10643 3451
rect 17969 3417 18003 3451
rect 19717 3417 19751 3451
rect 21373 3417 21407 3451
rect 46489 3417 46523 3451
rect 9045 3349 9079 3383
rect 14197 3349 14231 3383
rect 17325 3349 17359 3383
rect 28365 3349 28399 3383
rect 32321 3349 32355 3383
rect 45109 3349 45143 3383
rect 10701 3145 10735 3179
rect 47685 3145 47719 3179
rect 1869 3077 1903 3111
rect 4169 3077 4203 3111
rect 8033 3077 8067 3111
rect 13645 3077 13679 3111
rect 17325 3077 17359 3111
rect 19625 3077 19659 3111
rect 38761 3077 38795 3111
rect 42625 3077 42659 3111
rect 1685 3009 1719 3043
rect 6561 3009 6595 3043
rect 7849 3009 7883 3043
rect 10609 3009 10643 3043
rect 12633 3009 12667 3043
rect 13461 3009 13495 3043
rect 17141 3009 17175 3043
rect 22017 3009 22051 3043
rect 25605 3009 25639 3043
rect 32137 3009 32171 3043
rect 38577 3009 38611 3043
rect 41705 3009 41739 3043
rect 44741 3009 44775 3043
rect 47593 3009 47627 3043
rect 2789 2941 2823 2975
rect 3985 2941 4019 2975
rect 4813 2941 4847 2975
rect 8493 2941 8527 2975
rect 13921 2941 13955 2975
rect 17601 2941 17635 2975
rect 19441 2941 19475 2975
rect 20637 2941 20671 2975
rect 22201 2941 22235 2975
rect 22569 2941 22603 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 27169 2941 27203 2975
rect 27445 2941 27479 2975
rect 32321 2941 32355 2975
rect 32597 2941 32631 2975
rect 39313 2941 39347 2975
rect 41061 2941 41095 2975
rect 42441 2941 42475 2975
rect 42901 2941 42935 2975
rect 44925 2941 44959 2975
rect 46581 2941 46615 2975
rect 6653 2805 6687 2839
rect 7389 2805 7423 2839
rect 41797 2805 41831 2839
rect 2421 2601 2455 2635
rect 19901 2601 19935 2635
rect 47777 2601 47811 2635
rect 1777 2533 1811 2567
rect 4261 2465 4295 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 6837 2465 6871 2499
rect 8953 2465 8987 2499
rect 9137 2465 9171 2499
rect 9413 2465 9447 2499
rect 24685 2465 24719 2499
rect 27169 2465 27203 2499
rect 27353 2465 27387 2499
rect 28549 2465 28583 2499
rect 42441 2465 42475 2499
rect 42625 2465 42659 2499
rect 45017 2465 45051 2499
rect 45201 2465 45235 2499
rect 45569 2465 45603 2499
rect 3249 2397 3283 2431
rect 3801 2397 3835 2431
rect 24409 2397 24443 2431
rect 3985 2329 4019 2363
rect 44281 2329 44315 2363
<< metal1 >>
rect 38654 47404 38660 47456
rect 38712 47444 38718 47456
rect 39942 47444 39948 47456
rect 38712 47416 39948 47444
rect 38712 47404 38718 47416
rect 39942 47404 39948 47416
rect 40000 47404 40006 47456
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 2958 47132 2964 47184
rect 3016 47172 3022 47184
rect 4893 47175 4951 47181
rect 4893 47172 4905 47175
rect 3016 47144 4905 47172
rect 3016 47132 3022 47144
rect 4893 47141 4905 47144
rect 4939 47141 4951 47175
rect 4893 47135 4951 47141
rect 27614 47132 27620 47184
rect 27672 47172 27678 47184
rect 27801 47175 27859 47181
rect 27801 47172 27813 47175
rect 27672 47144 27813 47172
rect 27672 47132 27678 47144
rect 27801 47141 27813 47144
rect 27847 47141 27859 47175
rect 27801 47135 27859 47141
rect 45186 47132 45192 47184
rect 45244 47172 45250 47184
rect 47029 47175 47087 47181
rect 47029 47172 47041 47175
rect 45244 47144 47041 47172
rect 45244 47132 45250 47144
rect 47029 47141 47041 47144
rect 47075 47141 47087 47175
rect 47029 47135 47087 47141
rect 14 47064 20 47116
rect 72 47104 78 47116
rect 1397 47107 1455 47113
rect 1397 47104 1409 47107
rect 72 47076 1409 47104
rect 72 47064 78 47076
rect 1397 47073 1409 47076
rect 1443 47073 1455 47107
rect 11514 47104 11520 47116
rect 1397 47067 1455 47073
rect 2792 47076 11520 47104
rect 1673 47039 1731 47045
rect 1673 47005 1685 47039
rect 1719 47036 1731 47039
rect 2682 47036 2688 47048
rect 1719 47008 2688 47036
rect 1719 47005 1731 47008
rect 1673 46999 1731 47005
rect 2682 46996 2688 47008
rect 2740 46996 2746 47048
rect 2792 47045 2820 47076
rect 11514 47064 11520 47076
rect 11572 47064 11578 47116
rect 28810 47064 28816 47116
rect 28868 47104 28874 47116
rect 46842 47104 46848 47116
rect 28868 47076 46848 47104
rect 28868 47064 28874 47076
rect 46842 47064 46848 47076
rect 46900 47064 46906 47116
rect 2777 47039 2835 47045
rect 2777 47005 2789 47039
rect 2823 47005 2835 47039
rect 4246 47036 4252 47048
rect 4207 47008 4252 47036
rect 2777 46999 2835 47005
rect 4246 46996 4252 47008
rect 4304 46996 4310 47048
rect 5534 47036 5540 47048
rect 5495 47008 5540 47036
rect 5534 46996 5540 47008
rect 5592 46996 5598 47048
rect 8386 46996 8392 47048
rect 8444 47036 8450 47048
rect 9125 47039 9183 47045
rect 9125 47036 9137 47039
rect 8444 47008 9137 47036
rect 8444 46996 8450 47008
rect 9125 47005 9137 47008
rect 9171 47005 9183 47039
rect 12710 47036 12716 47048
rect 12671 47008 12716 47036
rect 9125 46999 9183 47005
rect 12710 46996 12716 47008
rect 12768 46996 12774 47048
rect 13170 46996 13176 47048
rect 13228 47036 13234 47048
rect 13449 47039 13507 47045
rect 13449 47036 13461 47039
rect 13228 47008 13461 47036
rect 13228 46996 13234 47008
rect 13449 47005 13461 47008
rect 13495 47005 13507 47039
rect 13449 46999 13507 47005
rect 14182 46996 14188 47048
rect 14240 47036 14246 47048
rect 14461 47039 14519 47045
rect 14461 47036 14473 47039
rect 14240 47008 14473 47036
rect 14240 46996 14246 47008
rect 14461 47005 14473 47008
rect 14507 47005 14519 47039
rect 15654 47036 15660 47048
rect 15615 47008 15660 47036
rect 14461 46999 14519 47005
rect 15654 46996 15660 47008
rect 15712 46996 15718 47048
rect 24854 47036 24860 47048
rect 24815 47008 24860 47036
rect 24854 46996 24860 47008
rect 24912 46996 24918 47048
rect 25498 47036 25504 47048
rect 25459 47008 25504 47036
rect 25498 46996 25504 47008
rect 25556 46996 25562 47048
rect 26418 47036 26424 47048
rect 26379 47008 26424 47036
rect 26418 46996 26424 47008
rect 26476 46996 26482 47048
rect 27982 47036 27988 47048
rect 27943 47008 27988 47036
rect 27982 46996 27988 47008
rect 28040 46996 28046 47048
rect 29730 46996 29736 47048
rect 29788 47036 29794 47048
rect 30101 47039 30159 47045
rect 30101 47036 30113 47039
rect 29788 47008 30113 47036
rect 29788 46996 29794 47008
rect 30101 47005 30113 47008
rect 30147 47005 30159 47039
rect 30101 46999 30159 47005
rect 32766 46996 32772 47048
rect 32824 47036 32830 47048
rect 33045 47039 33103 47045
rect 33045 47036 33057 47039
rect 32824 47008 33057 47036
rect 32824 46996 32830 47008
rect 33045 47005 33057 47008
rect 33091 47005 33103 47039
rect 33045 46999 33103 47005
rect 36081 47039 36139 47045
rect 36081 47005 36093 47039
rect 36127 47036 36139 47039
rect 37274 47036 37280 47048
rect 36127 47008 37280 47036
rect 36127 47005 36139 47008
rect 36081 46999 36139 47005
rect 37274 46996 37280 47008
rect 37332 46996 37338 47048
rect 46382 47036 46388 47048
rect 46343 47008 46388 47036
rect 46382 46996 46388 47008
rect 46440 46996 46446 47048
rect 47118 46996 47124 47048
rect 47176 47036 47182 47048
rect 47581 47039 47639 47045
rect 47581 47036 47593 47039
rect 47176 47008 47593 47036
rect 47176 46996 47182 47008
rect 47581 47005 47593 47008
rect 47627 47005 47639 47039
rect 47581 46999 47639 47005
rect 2866 46968 2872 46980
rect 2827 46940 2872 46968
rect 2866 46928 2872 46940
rect 2924 46928 2930 46980
rect 46566 46928 46572 46980
rect 46624 46968 46630 46980
rect 47673 46971 47731 46977
rect 47673 46968 47685 46971
rect 46624 46940 47685 46968
rect 46624 46928 46630 46940
rect 47673 46937 47685 46940
rect 47719 46937 47731 46971
rect 47673 46931 47731 46937
rect 8938 46900 8944 46912
rect 8899 46872 8944 46900
rect 8938 46860 8944 46872
rect 8996 46860 9002 46912
rect 40586 46860 40592 46912
rect 40644 46900 40650 46912
rect 41414 46900 41420 46912
rect 40644 46872 41420 46900
rect 40644 46860 40650 46872
rect 41414 46860 41420 46872
rect 41472 46860 41478 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 2590 46656 2596 46708
rect 2648 46696 2654 46708
rect 3050 46696 3056 46708
rect 2648 46668 3056 46696
rect 2648 46656 2654 46668
rect 3050 46656 3056 46668
rect 3108 46656 3114 46708
rect 1857 46631 1915 46637
rect 1857 46597 1869 46631
rect 1903 46628 1915 46631
rect 3878 46628 3884 46640
rect 1903 46600 3884 46628
rect 1903 46597 1915 46600
rect 1857 46591 1915 46597
rect 3878 46588 3884 46600
rect 3936 46588 3942 46640
rect 4246 46628 4252 46640
rect 3988 46600 4252 46628
rect 3988 46569 4016 46600
rect 4246 46588 4252 46600
rect 4304 46588 4310 46640
rect 12710 46628 12716 46640
rect 11900 46600 12716 46628
rect 11900 46569 11928 46600
rect 12710 46588 12716 46600
rect 12768 46588 12774 46640
rect 25498 46628 25504 46640
rect 24596 46600 25504 46628
rect 3973 46563 4031 46569
rect 3973 46529 3985 46563
rect 4019 46529 4031 46563
rect 3973 46523 4031 46529
rect 11885 46563 11943 46569
rect 11885 46529 11897 46563
rect 11931 46529 11943 46563
rect 14182 46560 14188 46572
rect 14143 46532 14188 46560
rect 11885 46523 11943 46529
rect 14182 46520 14188 46532
rect 14240 46520 14246 46572
rect 24596 46569 24624 46600
rect 25498 46588 25504 46600
rect 25556 46588 25562 46640
rect 46382 46628 46388 46640
rect 45204 46600 46388 46628
rect 24581 46563 24639 46569
rect 24581 46529 24593 46563
rect 24627 46529 24639 46563
rect 24581 46523 24639 46529
rect 26418 46520 26424 46572
rect 26476 46560 26482 46572
rect 26973 46563 27031 46569
rect 26973 46560 26985 46563
rect 26476 46532 26985 46560
rect 26476 46520 26482 46532
rect 26973 46529 26985 46532
rect 27019 46529 27031 46563
rect 29730 46560 29736 46572
rect 29691 46532 29736 46560
rect 26973 46523 27031 46529
rect 29730 46520 29736 46532
rect 29788 46520 29794 46572
rect 32766 46560 32772 46572
rect 32727 46532 32772 46560
rect 32766 46520 32772 46532
rect 32824 46520 32830 46572
rect 35802 46560 35808 46572
rect 35763 46532 35808 46560
rect 35802 46520 35808 46532
rect 35860 46520 35866 46572
rect 37274 46560 37280 46572
rect 37235 46532 37280 46560
rect 37274 46520 37280 46532
rect 37332 46520 37338 46572
rect 45204 46569 45232 46600
rect 46382 46588 46388 46600
rect 46440 46588 46446 46640
rect 45189 46563 45247 46569
rect 45189 46529 45201 46563
rect 45235 46529 45247 46563
rect 45189 46523 45247 46529
rect 47210 46520 47216 46572
rect 47268 46560 47274 46572
rect 47581 46563 47639 46569
rect 47581 46560 47593 46563
rect 47268 46532 47593 46560
rect 47268 46520 47274 46532
rect 47581 46529 47593 46532
rect 47627 46529 47639 46563
rect 47581 46523 47639 46529
rect 1673 46495 1731 46501
rect 1673 46461 1685 46495
rect 1719 46492 1731 46495
rect 2130 46492 2136 46504
rect 1719 46464 1808 46492
rect 2091 46464 2136 46492
rect 1719 46461 1731 46464
rect 1673 46455 1731 46461
rect 1780 46436 1808 46464
rect 2130 46452 2136 46464
rect 2188 46452 2194 46504
rect 4157 46495 4215 46501
rect 4157 46461 4169 46495
rect 4203 46461 4215 46495
rect 4614 46492 4620 46504
rect 4575 46464 4620 46492
rect 4157 46455 4215 46461
rect 1762 46384 1768 46436
rect 1820 46384 1826 46436
rect 4062 46384 4068 46436
rect 4120 46424 4126 46436
rect 4172 46424 4200 46455
rect 4614 46452 4620 46464
rect 4672 46452 4678 46504
rect 12069 46495 12127 46501
rect 12069 46461 12081 46495
rect 12115 46492 12127 46495
rect 12618 46492 12624 46504
rect 12115 46464 12624 46492
rect 12115 46461 12127 46464
rect 12069 46455 12127 46461
rect 12618 46452 12624 46464
rect 12676 46452 12682 46504
rect 12894 46492 12900 46504
rect 12855 46464 12900 46492
rect 12894 46452 12900 46464
rect 12952 46452 12958 46504
rect 14369 46495 14427 46501
rect 14369 46461 14381 46495
rect 14415 46492 14427 46495
rect 14458 46492 14464 46504
rect 14415 46464 14464 46492
rect 14415 46461 14427 46464
rect 14369 46455 14427 46461
rect 14458 46452 14464 46464
rect 14516 46452 14522 46504
rect 14826 46492 14832 46504
rect 14787 46464 14832 46492
rect 14826 46452 14832 46464
rect 14884 46452 14890 46504
rect 22278 46492 22284 46504
rect 22239 46464 22284 46492
rect 22278 46452 22284 46464
rect 22336 46452 22342 46504
rect 22465 46495 22523 46501
rect 22465 46461 22477 46495
rect 22511 46492 22523 46495
rect 22922 46492 22928 46504
rect 22511 46464 22928 46492
rect 22511 46461 22523 46464
rect 22465 46455 22523 46461
rect 22922 46452 22928 46464
rect 22980 46452 22986 46504
rect 23198 46492 23204 46504
rect 23159 46464 23204 46492
rect 23198 46452 23204 46464
rect 23256 46452 23262 46504
rect 24765 46495 24823 46501
rect 24765 46461 24777 46495
rect 24811 46492 24823 46495
rect 25314 46492 25320 46504
rect 24811 46464 25320 46492
rect 24811 46461 24823 46464
rect 24765 46455 24823 46461
rect 25314 46452 25320 46464
rect 25372 46452 25378 46504
rect 25774 46492 25780 46504
rect 25735 46464 25780 46492
rect 25774 46452 25780 46464
rect 25832 46452 25838 46504
rect 26234 46452 26240 46504
rect 26292 46492 26298 46504
rect 27157 46495 27215 46501
rect 27157 46492 27169 46495
rect 26292 46464 27169 46492
rect 26292 46452 26298 46464
rect 27157 46461 27169 46464
rect 27203 46461 27215 46495
rect 27157 46455 27215 46461
rect 27617 46495 27675 46501
rect 27617 46461 27629 46495
rect 27663 46461 27675 46495
rect 29914 46492 29920 46504
rect 29875 46464 29920 46492
rect 27617 46455 27675 46461
rect 4120 46396 4200 46424
rect 4120 46384 4126 46396
rect 9582 46384 9588 46436
rect 9640 46424 9646 46436
rect 17218 46424 17224 46436
rect 9640 46396 17224 46424
rect 9640 46384 9646 46396
rect 17218 46384 17224 46396
rect 17276 46384 17282 46436
rect 27062 46384 27068 46436
rect 27120 46424 27126 46436
rect 27632 46424 27660 46455
rect 29914 46452 29920 46464
rect 29972 46452 29978 46504
rect 30282 46452 30288 46504
rect 30340 46492 30346 46504
rect 30377 46495 30435 46501
rect 30377 46492 30389 46495
rect 30340 46464 30389 46492
rect 30340 46452 30346 46464
rect 30377 46461 30389 46464
rect 30423 46461 30435 46495
rect 32950 46492 32956 46504
rect 32911 46464 32956 46492
rect 30377 46455 30435 46461
rect 32950 46452 32956 46464
rect 33008 46452 33014 46504
rect 33502 46492 33508 46504
rect 33463 46464 33508 46492
rect 33502 46452 33508 46464
rect 33560 46452 33566 46504
rect 37458 46492 37464 46504
rect 37419 46464 37464 46492
rect 37458 46452 37464 46464
rect 37516 46452 37522 46504
rect 37737 46495 37795 46501
rect 37737 46461 37749 46495
rect 37783 46461 37795 46495
rect 37737 46455 37795 46461
rect 45373 46495 45431 46501
rect 45373 46461 45385 46495
rect 45419 46492 45431 46495
rect 46566 46492 46572 46504
rect 45419 46464 46572 46492
rect 45419 46461 45431 46464
rect 45373 46455 45431 46461
rect 27120 46396 27660 46424
rect 27120 46384 27126 46396
rect 35710 46384 35716 46436
rect 35768 46424 35774 46436
rect 36633 46427 36691 46433
rect 36633 46424 36645 46427
rect 35768 46396 36645 46424
rect 35768 46384 35774 46396
rect 36633 46393 36645 46396
rect 36679 46393 36691 46427
rect 36633 46387 36691 46393
rect 36722 46384 36728 46436
rect 36780 46424 36786 46436
rect 37752 46424 37780 46455
rect 46566 46452 46572 46464
rect 46624 46452 46630 46504
rect 46750 46492 46756 46504
rect 46711 46464 46756 46492
rect 46750 46452 46756 46464
rect 46808 46452 46814 46504
rect 36780 46396 37780 46424
rect 36780 46384 36786 46396
rect 10870 46316 10876 46368
rect 10928 46356 10934 46368
rect 10965 46359 11023 46365
rect 10965 46356 10977 46359
rect 10928 46328 10977 46356
rect 10928 46316 10934 46328
rect 10965 46325 10977 46328
rect 11011 46325 11023 46359
rect 10965 46319 11023 46325
rect 35894 46316 35900 46368
rect 35952 46356 35958 46368
rect 35952 46328 35997 46356
rect 35952 46316 35958 46328
rect 41598 46316 41604 46368
rect 41656 46356 41662 46368
rect 41785 46359 41843 46365
rect 41785 46356 41797 46359
rect 41656 46328 41797 46356
rect 41656 46316 41662 46328
rect 41785 46325 41797 46328
rect 41831 46325 41843 46359
rect 41785 46319 41843 46325
rect 45646 46316 45652 46368
rect 45704 46356 45710 46368
rect 47673 46359 47731 46365
rect 47673 46356 47685 46359
rect 45704 46328 47685 46356
rect 45704 46316 45710 46328
rect 47673 46325 47685 46328
rect 47719 46325 47731 46359
rect 47673 46319 47731 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 4062 46112 4068 46164
rect 4120 46152 4126 46164
rect 4157 46155 4215 46161
rect 4157 46152 4169 46155
rect 4120 46124 4169 46152
rect 4120 46112 4126 46124
rect 4157 46121 4169 46124
rect 4203 46121 4215 46155
rect 14458 46152 14464 46164
rect 14419 46124 14464 46152
rect 4157 46115 4215 46121
rect 14458 46112 14464 46124
rect 14516 46112 14522 46164
rect 22278 46112 22284 46164
rect 22336 46152 22342 46164
rect 23017 46155 23075 46161
rect 23017 46152 23029 46155
rect 22336 46124 23029 46152
rect 22336 46112 22342 46124
rect 23017 46121 23029 46124
rect 23063 46121 23075 46155
rect 23017 46115 23075 46121
rect 32861 46155 32919 46161
rect 32861 46121 32873 46155
rect 32907 46152 32919 46155
rect 32950 46152 32956 46164
rect 32907 46124 32956 46152
rect 32907 46121 32919 46124
rect 32861 46115 32919 46121
rect 32950 46112 32956 46124
rect 33008 46112 33014 46164
rect 47210 46152 47216 46164
rect 35866 46124 47216 46152
rect 10962 46044 10968 46096
rect 11020 46044 11026 46096
rect 15470 46044 15476 46096
rect 15528 46084 15534 46096
rect 15528 46056 15884 46084
rect 15528 46044 15534 46056
rect 2774 46016 2780 46028
rect 2735 45988 2780 46016
rect 2774 45976 2780 45988
rect 2832 45976 2838 46028
rect 5261 46019 5319 46025
rect 5261 45985 5273 46019
rect 5307 46016 5319 46019
rect 5534 46016 5540 46028
rect 5307 45988 5540 46016
rect 5307 45985 5319 45988
rect 5261 45979 5319 45985
rect 5534 45976 5540 45988
rect 5592 45976 5598 46028
rect 5810 46016 5816 46028
rect 5771 45988 5816 46016
rect 5810 45976 5816 45988
rect 5868 45976 5874 46028
rect 9582 46016 9588 46028
rect 9543 45988 9588 46016
rect 9582 45976 9588 45988
rect 9640 45976 9646 46028
rect 10870 46016 10876 46028
rect 10831 45988 10876 46016
rect 10870 45976 10876 45988
rect 10928 45976 10934 46028
rect 10980 46016 11008 46044
rect 11333 46019 11391 46025
rect 11333 46016 11345 46019
rect 10980 45988 11345 46016
rect 11333 45985 11345 45988
rect 11379 45985 11391 46019
rect 11333 45979 11391 45985
rect 15381 46019 15439 46025
rect 15381 45985 15393 46019
rect 15427 46016 15439 46019
rect 15654 46016 15660 46028
rect 15427 45988 15660 46016
rect 15427 45985 15439 45988
rect 15381 45979 15439 45985
rect 15654 45976 15660 45988
rect 15712 45976 15718 46028
rect 15856 46025 15884 46056
rect 15841 46019 15899 46025
rect 15841 45985 15853 46019
rect 15887 45985 15899 46019
rect 15841 45979 15899 45985
rect 17218 45976 17224 46028
rect 17276 46016 17282 46028
rect 35866 46016 35894 46124
rect 47210 46112 47216 46124
rect 47268 46112 47274 46164
rect 17276 45988 35894 46016
rect 17276 45976 17282 45988
rect 36078 45976 36084 46028
rect 36136 46016 36142 46028
rect 36173 46019 36231 46025
rect 36173 46016 36185 46019
rect 36136 45988 36185 46016
rect 36136 45976 36142 45988
rect 36173 45985 36185 45988
rect 36219 45985 36231 46019
rect 41598 46016 41604 46028
rect 41559 45988 41604 46016
rect 36173 45979 36231 45985
rect 41598 45976 41604 45988
rect 41656 45976 41662 46028
rect 42058 46016 42064 46028
rect 42019 45988 42064 46016
rect 42058 45976 42064 45988
rect 42116 45976 42122 46028
rect 48133 46019 48191 46025
rect 48133 45985 48145 46019
rect 48179 46016 48191 46019
rect 48314 46016 48320 46028
rect 48179 45988 48320 46016
rect 48179 45985 48191 45988
rect 48133 45979 48191 45985
rect 48314 45976 48320 45988
rect 48372 45976 48378 46028
rect 1394 45948 1400 45960
rect 1355 45920 1400 45948
rect 1394 45908 1400 45920
rect 1452 45908 1458 45960
rect 4065 45951 4123 45957
rect 4065 45917 4077 45951
rect 4111 45917 4123 45951
rect 9214 45948 9220 45960
rect 9175 45920 9220 45948
rect 4065 45911 4123 45917
rect 1581 45883 1639 45889
rect 1581 45849 1593 45883
rect 1627 45880 1639 45883
rect 3142 45880 3148 45892
rect 1627 45852 3148 45880
rect 1627 45849 1639 45852
rect 1581 45843 1639 45849
rect 3142 45840 3148 45852
rect 3200 45840 3206 45892
rect 4080 45824 4108 45911
rect 9214 45908 9220 45920
rect 9272 45908 9278 45960
rect 12526 45908 12532 45960
rect 12584 45948 12590 45960
rect 13173 45951 13231 45957
rect 13173 45948 13185 45951
rect 12584 45920 13185 45948
rect 12584 45908 12590 45920
rect 13173 45917 13185 45920
rect 13219 45917 13231 45951
rect 13173 45911 13231 45917
rect 14369 45951 14427 45957
rect 14369 45917 14381 45951
rect 14415 45917 14427 45951
rect 24670 45948 24676 45960
rect 24631 45920 24676 45948
rect 14369 45911 14427 45917
rect 5445 45883 5503 45889
rect 5445 45849 5457 45883
rect 5491 45880 5503 45883
rect 5534 45880 5540 45892
rect 5491 45852 5540 45880
rect 5491 45849 5503 45852
rect 5445 45843 5503 45849
rect 5534 45840 5540 45852
rect 5592 45840 5598 45892
rect 11057 45883 11115 45889
rect 11057 45849 11069 45883
rect 11103 45880 11115 45883
rect 11606 45880 11612 45892
rect 11103 45852 11612 45880
rect 11103 45849 11115 45852
rect 11057 45843 11115 45849
rect 11606 45840 11612 45852
rect 11664 45840 11670 45892
rect 14384 45824 14412 45911
rect 24670 45908 24676 45920
rect 24728 45908 24734 45960
rect 26970 45948 26976 45960
rect 26931 45920 26976 45948
rect 26970 45908 26976 45920
rect 27028 45908 27034 45960
rect 28810 45948 28816 45960
rect 28771 45920 28816 45948
rect 28810 45908 28816 45920
rect 28868 45908 28874 45960
rect 29730 45948 29736 45960
rect 29691 45920 29736 45948
rect 29730 45908 29736 45920
rect 29788 45908 29794 45960
rect 32766 45948 32772 45960
rect 32727 45920 32772 45948
rect 32766 45908 32772 45920
rect 32824 45908 32830 45960
rect 35710 45948 35716 45960
rect 35671 45920 35716 45948
rect 35710 45908 35716 45920
rect 35768 45908 35774 45960
rect 38102 45908 38108 45960
rect 38160 45948 38166 45960
rect 38289 45951 38347 45957
rect 38289 45948 38301 45951
rect 38160 45920 38301 45948
rect 38160 45908 38166 45920
rect 38289 45917 38301 45920
rect 38335 45917 38347 45951
rect 38289 45911 38347 45917
rect 45833 45951 45891 45957
rect 45833 45917 45845 45951
rect 45879 45948 45891 45951
rect 46293 45951 46351 45957
rect 46293 45948 46305 45951
rect 45879 45920 46305 45948
rect 45879 45917 45891 45920
rect 45833 45911 45891 45917
rect 46293 45917 46305 45920
rect 46339 45917 46351 45951
rect 46293 45911 46351 45917
rect 15562 45880 15568 45892
rect 15523 45852 15568 45880
rect 15562 45840 15568 45852
rect 15620 45840 15626 45892
rect 24854 45880 24860 45892
rect 24815 45852 24860 45880
rect 24854 45840 24860 45852
rect 24912 45840 24918 45892
rect 25130 45840 25136 45892
rect 25188 45880 25194 45892
rect 26513 45883 26571 45889
rect 26513 45880 26525 45883
rect 25188 45852 26525 45880
rect 25188 45840 25194 45852
rect 26513 45849 26525 45852
rect 26559 45849 26571 45883
rect 27154 45880 27160 45892
rect 27115 45852 27160 45880
rect 26513 45843 26571 45849
rect 27154 45840 27160 45852
rect 27212 45840 27218 45892
rect 35894 45840 35900 45892
rect 35952 45880 35958 45892
rect 41782 45880 41788 45892
rect 35952 45852 35997 45880
rect 41743 45852 41788 45880
rect 35952 45840 35958 45852
rect 41782 45840 41788 45852
rect 41840 45840 41846 45892
rect 46477 45883 46535 45889
rect 46477 45849 46489 45883
rect 46523 45880 46535 45883
rect 47670 45880 47676 45892
rect 46523 45852 47676 45880
rect 46523 45849 46535 45852
rect 46477 45843 46535 45849
rect 47670 45840 47676 45852
rect 47728 45840 47734 45892
rect 4062 45812 4068 45824
rect 3975 45784 4068 45812
rect 4062 45772 4068 45784
rect 4120 45812 4126 45824
rect 10778 45812 10784 45824
rect 4120 45784 10784 45812
rect 4120 45772 4126 45784
rect 10778 45772 10784 45784
rect 10836 45772 10842 45824
rect 13265 45815 13323 45821
rect 13265 45781 13277 45815
rect 13311 45812 13323 45815
rect 13354 45812 13360 45824
rect 13311 45784 13360 45812
rect 13311 45781 13323 45784
rect 13265 45775 13323 45781
rect 13354 45772 13360 45784
rect 13412 45772 13418 45824
rect 14366 45812 14372 45824
rect 14279 45784 14372 45812
rect 14366 45772 14372 45784
rect 14424 45812 14430 45824
rect 35802 45812 35808 45824
rect 14424 45784 35808 45812
rect 14424 45772 14430 45784
rect 35802 45772 35808 45784
rect 35860 45772 35866 45824
rect 40678 45772 40684 45824
rect 40736 45812 40742 45824
rect 47118 45812 47124 45824
rect 40736 45784 47124 45812
rect 40736 45772 40742 45784
rect 47118 45772 47124 45784
rect 47176 45772 47182 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 11606 45608 11612 45620
rect 11567 45580 11612 45608
rect 11606 45568 11612 45580
rect 11664 45568 11670 45620
rect 13188 45580 13492 45608
rect 1670 45540 1676 45552
rect 1631 45512 1676 45540
rect 1670 45500 1676 45512
rect 1728 45500 1734 45552
rect 2501 45543 2559 45549
rect 2501 45509 2513 45543
rect 2547 45540 2559 45543
rect 2866 45540 2872 45552
rect 2547 45512 2872 45540
rect 2547 45509 2559 45512
rect 2501 45503 2559 45509
rect 2866 45500 2872 45512
rect 2924 45500 2930 45552
rect 5534 45540 5540 45552
rect 5495 45512 5540 45540
rect 5534 45500 5540 45512
rect 5592 45500 5598 45552
rect 9582 45540 9588 45552
rect 6886 45512 9588 45540
rect 5442 45472 5448 45484
rect 5403 45444 5448 45472
rect 5442 45432 5448 45444
rect 5500 45472 5506 45484
rect 6886 45472 6914 45512
rect 9582 45500 9588 45512
rect 9640 45500 9646 45552
rect 12618 45540 12624 45552
rect 12579 45512 12624 45540
rect 12618 45500 12624 45512
rect 12676 45500 12682 45552
rect 13188 45540 13216 45580
rect 13354 45540 13360 45552
rect 13004 45512 13216 45540
rect 13315 45512 13360 45540
rect 8386 45472 8392 45484
rect 5500 45444 6914 45472
rect 8347 45444 8392 45472
rect 5500 45432 5506 45444
rect 8386 45432 8392 45444
rect 8444 45432 8450 45484
rect 8573 45475 8631 45481
rect 8573 45441 8585 45475
rect 8619 45472 8631 45475
rect 9125 45475 9183 45481
rect 9125 45472 9137 45475
rect 8619 45444 9137 45472
rect 8619 45441 8631 45444
rect 8573 45435 8631 45441
rect 9125 45441 9137 45444
rect 9171 45472 9183 45475
rect 9214 45472 9220 45484
rect 9171 45444 9220 45472
rect 9171 45441 9183 45444
rect 9125 45435 9183 45441
rect 9214 45432 9220 45444
rect 9272 45472 9278 45484
rect 10321 45475 10379 45481
rect 10321 45472 10333 45475
rect 9272 45444 10333 45472
rect 9272 45432 9278 45444
rect 10321 45441 10333 45444
rect 10367 45441 10379 45475
rect 11514 45472 11520 45484
rect 11427 45444 11520 45472
rect 10321 45435 10379 45441
rect 11514 45432 11520 45444
rect 11572 45432 11578 45484
rect 12526 45472 12532 45484
rect 12487 45444 12532 45472
rect 12526 45432 12532 45444
rect 12584 45432 12590 45484
rect 2317 45407 2375 45413
rect 2317 45373 2329 45407
rect 2363 45404 2375 45407
rect 2958 45404 2964 45416
rect 2363 45376 2964 45404
rect 2363 45373 2375 45376
rect 2317 45367 2375 45373
rect 2958 45364 2964 45376
rect 3016 45364 3022 45416
rect 3050 45364 3056 45416
rect 3108 45404 3114 45416
rect 9398 45404 9404 45416
rect 3108 45376 3153 45404
rect 9359 45376 9404 45404
rect 3108 45364 3114 45376
rect 9398 45364 9404 45376
rect 9456 45364 9462 45416
rect 10778 45364 10784 45416
rect 10836 45404 10842 45416
rect 10873 45407 10931 45413
rect 10873 45404 10885 45407
rect 10836 45376 10885 45404
rect 10836 45364 10842 45376
rect 10873 45373 10885 45376
rect 10919 45373 10931 45407
rect 11532 45404 11560 45432
rect 13004 45404 13032 45512
rect 13354 45500 13360 45512
rect 13412 45500 13418 45552
rect 13464 45540 13492 45580
rect 15562 45568 15568 45620
rect 15620 45608 15626 45620
rect 15657 45611 15715 45617
rect 15657 45608 15669 45611
rect 15620 45580 15669 45608
rect 15620 45568 15626 45580
rect 15657 45577 15669 45580
rect 15703 45577 15715 45611
rect 22922 45608 22928 45620
rect 22883 45580 22928 45608
rect 15657 45571 15715 45577
rect 22922 45568 22928 45580
rect 22980 45568 22986 45620
rect 32766 45568 32772 45620
rect 32824 45608 32830 45620
rect 40678 45608 40684 45620
rect 32824 45580 40684 45608
rect 32824 45568 32830 45580
rect 40678 45568 40684 45580
rect 40736 45568 40742 45620
rect 18506 45540 18512 45552
rect 13464 45512 18512 45540
rect 18506 45500 18512 45512
rect 18564 45500 18570 45552
rect 24673 45543 24731 45549
rect 24673 45509 24685 45543
rect 24719 45540 24731 45543
rect 24854 45540 24860 45552
rect 24719 45512 24860 45540
rect 24719 45509 24731 45512
rect 24673 45503 24731 45509
rect 24854 45500 24860 45512
rect 24912 45500 24918 45552
rect 25314 45540 25320 45552
rect 25275 45512 25320 45540
rect 25314 45500 25320 45512
rect 25372 45500 25378 45552
rect 29730 45540 29736 45552
rect 25424 45512 27384 45540
rect 13170 45472 13176 45484
rect 13131 45444 13176 45472
rect 13170 45432 13176 45444
rect 13228 45432 13234 45484
rect 15562 45472 15568 45484
rect 15475 45444 15568 45472
rect 15562 45432 15568 45444
rect 15620 45472 15626 45484
rect 22830 45472 22836 45484
rect 15620 45444 22094 45472
rect 22791 45444 22836 45472
rect 15620 45432 15626 45444
rect 14274 45404 14280 45416
rect 11532 45376 13032 45404
rect 14235 45376 14280 45404
rect 10873 45367 10931 45373
rect 1857 45339 1915 45345
rect 1857 45305 1869 45339
rect 1903 45336 1915 45339
rect 8386 45336 8392 45348
rect 1903 45308 8392 45336
rect 1903 45305 1915 45308
rect 1857 45299 1915 45305
rect 8386 45296 8392 45308
rect 8444 45296 8450 45348
rect 10888 45336 10916 45367
rect 14274 45364 14280 45376
rect 14332 45364 14338 45416
rect 22066 45404 22094 45444
rect 22830 45432 22836 45444
rect 22888 45432 22894 45484
rect 24486 45432 24492 45484
rect 24544 45472 24550 45484
rect 24581 45475 24639 45481
rect 24581 45472 24593 45475
rect 24544 45444 24593 45472
rect 24544 45432 24550 45444
rect 24581 45441 24593 45444
rect 24627 45472 24639 45475
rect 25225 45475 25283 45481
rect 25225 45472 25237 45475
rect 24627 45444 25237 45472
rect 24627 45441 24639 45444
rect 24581 45435 24639 45441
rect 25225 45441 25237 45444
rect 25271 45441 25283 45475
rect 25225 45435 25283 45441
rect 25424 45404 25452 45512
rect 26053 45475 26111 45481
rect 26053 45441 26065 45475
rect 26099 45441 26111 45475
rect 26053 45435 26111 45441
rect 26145 45475 26203 45481
rect 26145 45441 26157 45475
rect 26191 45472 26203 45475
rect 26234 45472 26240 45484
rect 26191 45444 26240 45472
rect 26191 45441 26203 45444
rect 26145 45435 26203 45441
rect 22066 45376 25452 45404
rect 26068 45348 26096 45435
rect 26234 45432 26240 45444
rect 26292 45432 26298 45484
rect 26970 45432 26976 45484
rect 27028 45472 27034 45484
rect 27249 45475 27307 45481
rect 27249 45472 27261 45475
rect 27028 45444 27261 45472
rect 27028 45432 27034 45444
rect 27249 45441 27261 45444
rect 27295 45441 27307 45475
rect 27249 45435 27307 45441
rect 26050 45336 26056 45348
rect 10888 45308 12434 45336
rect 12406 45268 12434 45308
rect 14200 45308 26056 45336
rect 14200 45268 14228 45308
rect 26050 45296 26056 45308
rect 26108 45296 26114 45348
rect 27356 45336 27384 45512
rect 28644 45512 29736 45540
rect 28644 45481 28672 45512
rect 29730 45500 29736 45512
rect 29788 45500 29794 45552
rect 39942 45540 39948 45552
rect 39903 45512 39948 45540
rect 39942 45500 39948 45512
rect 40000 45500 40006 45552
rect 45373 45543 45431 45549
rect 45373 45509 45385 45543
rect 45419 45540 45431 45543
rect 45646 45540 45652 45552
rect 45419 45512 45652 45540
rect 45419 45509 45431 45512
rect 45373 45503 45431 45509
rect 45646 45500 45652 45512
rect 45704 45500 45710 45552
rect 47670 45540 47676 45552
rect 47631 45512 47676 45540
rect 47670 45500 47676 45512
rect 47728 45500 47734 45552
rect 28629 45475 28687 45481
rect 28629 45441 28641 45475
rect 28675 45441 28687 45475
rect 28629 45435 28687 45441
rect 35921 45475 35979 45481
rect 35921 45441 35933 45475
rect 35967 45472 35979 45475
rect 36078 45472 36084 45484
rect 35967 45444 36084 45472
rect 35967 45441 35979 45444
rect 35921 45435 35979 45441
rect 36078 45432 36084 45444
rect 36136 45432 36142 45484
rect 38102 45472 38108 45484
rect 38063 45444 38108 45472
rect 38102 45432 38108 45444
rect 38160 45432 38166 45484
rect 45186 45472 45192 45484
rect 45147 45444 45192 45472
rect 45186 45432 45192 45444
rect 45244 45432 45250 45484
rect 47302 45432 47308 45484
rect 47360 45472 47366 45484
rect 47581 45475 47639 45481
rect 47581 45472 47593 45475
rect 47360 45444 47593 45472
rect 47360 45432 47366 45444
rect 47581 45441 47593 45444
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 27430 45364 27436 45416
rect 27488 45404 27494 45416
rect 28813 45407 28871 45413
rect 28813 45404 28825 45407
rect 27488 45376 28825 45404
rect 27488 45364 27494 45376
rect 28813 45373 28825 45376
rect 28859 45373 28871 45407
rect 30282 45404 30288 45416
rect 30243 45376 30288 45404
rect 28813 45367 28871 45373
rect 30282 45364 30288 45376
rect 30340 45364 30346 45416
rect 38010 45404 38016 45416
rect 35866 45376 38016 45404
rect 35866 45336 35894 45376
rect 38010 45364 38016 45376
rect 38068 45364 38074 45416
rect 38286 45404 38292 45416
rect 38247 45376 38292 45404
rect 38286 45364 38292 45376
rect 38344 45364 38350 45416
rect 46842 45404 46848 45416
rect 46803 45376 46848 45404
rect 46842 45364 46848 45376
rect 46900 45364 46906 45416
rect 27356 45308 35894 45336
rect 35989 45339 36047 45345
rect 35989 45305 36001 45339
rect 36035 45336 36047 45339
rect 37458 45336 37464 45348
rect 36035 45308 37464 45336
rect 36035 45305 36047 45308
rect 35989 45299 36047 45305
rect 37458 45296 37464 45308
rect 37516 45296 37522 45348
rect 12406 45240 14228 45268
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 1394 45024 1400 45076
rect 1452 45064 1458 45076
rect 1949 45067 2007 45073
rect 1949 45064 1961 45067
rect 1452 45036 1961 45064
rect 1452 45024 1458 45036
rect 1949 45033 1961 45036
rect 1995 45033 2007 45067
rect 3142 45064 3148 45076
rect 3103 45036 3148 45064
rect 1949 45027 2007 45033
rect 3142 45024 3148 45036
rect 3200 45024 3206 45076
rect 3878 45064 3884 45076
rect 3839 45036 3884 45064
rect 3878 45024 3884 45036
rect 3936 45024 3942 45076
rect 26789 45067 26847 45073
rect 26789 45033 26801 45067
rect 26835 45064 26847 45067
rect 27154 45064 27160 45076
rect 26835 45036 27160 45064
rect 26835 45033 26847 45036
rect 26789 45027 26847 45033
rect 27154 45024 27160 45036
rect 27212 45024 27218 45076
rect 27430 45064 27436 45076
rect 27391 45036 27436 45064
rect 27430 45024 27436 45036
rect 27488 45024 27494 45076
rect 29914 45024 29920 45076
rect 29972 45064 29978 45076
rect 30009 45067 30067 45073
rect 30009 45064 30021 45067
rect 29972 45036 30021 45064
rect 29972 45024 29978 45036
rect 30009 45033 30021 45036
rect 30055 45033 30067 45067
rect 30009 45027 30067 45033
rect 38197 45067 38255 45073
rect 38197 45033 38209 45067
rect 38243 45064 38255 45067
rect 38286 45064 38292 45076
rect 38243 45036 38292 45064
rect 38243 45033 38255 45036
rect 38197 45027 38255 45033
rect 38286 45024 38292 45036
rect 38344 45024 38350 45076
rect 41782 45064 41788 45076
rect 41743 45036 41788 45064
rect 41782 45024 41788 45036
rect 41840 45024 41846 45076
rect 1762 44956 1768 45008
rect 1820 44996 1826 45008
rect 2593 44999 2651 45005
rect 2593 44996 2605 44999
rect 1820 44968 2605 44996
rect 1820 44956 1826 44968
rect 2593 44965 2605 44968
rect 2639 44965 2651 44999
rect 2593 44959 2651 44965
rect 9398 44956 9404 45008
rect 9456 44996 9462 45008
rect 9456 44968 29960 44996
rect 9456 44956 9462 44968
rect 8202 44928 8208 44940
rect 6886 44900 8208 44928
rect 3050 44860 3056 44872
rect 3011 44832 3056 44860
rect 3050 44820 3056 44832
rect 3108 44820 3114 44872
rect 3789 44863 3847 44869
rect 3789 44829 3801 44863
rect 3835 44860 3847 44863
rect 6886 44860 6914 44900
rect 8202 44888 8208 44900
rect 8260 44928 8266 44940
rect 14366 44928 14372 44940
rect 8260 44900 14372 44928
rect 8260 44888 8266 44900
rect 14366 44888 14372 44900
rect 14424 44888 14430 44940
rect 29932 44872 29960 44968
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 9214 44860 9220 44872
rect 3835 44832 6914 44860
rect 9175 44832 9220 44860
rect 3835 44829 3847 44832
rect 3789 44823 3847 44829
rect 9214 44820 9220 44832
rect 9272 44820 9278 44872
rect 26694 44860 26700 44872
rect 26655 44832 26700 44860
rect 26694 44820 26700 44832
rect 26752 44860 26758 44872
rect 27341 44863 27399 44869
rect 27341 44860 27353 44863
rect 26752 44832 27353 44860
rect 26752 44820 26758 44832
rect 27341 44829 27353 44832
rect 27387 44829 27399 44863
rect 29914 44860 29920 44872
rect 29875 44832 29920 44860
rect 27341 44823 27399 44829
rect 29914 44820 29920 44832
rect 29972 44820 29978 44872
rect 38105 44863 38163 44869
rect 38105 44829 38117 44863
rect 38151 44860 38163 44863
rect 38286 44860 38292 44872
rect 38151 44832 38292 44860
rect 38151 44829 38163 44832
rect 38105 44823 38163 44829
rect 38286 44820 38292 44832
rect 38344 44820 38350 44872
rect 41693 44863 41751 44869
rect 41693 44829 41705 44863
rect 41739 44860 41751 44863
rect 41966 44860 41972 44872
rect 41739 44832 41972 44860
rect 41739 44829 41751 44832
rect 41693 44823 41751 44829
rect 41966 44820 41972 44832
rect 42024 44820 42030 44872
rect 45833 44863 45891 44869
rect 45833 44829 45845 44863
rect 45879 44860 45891 44863
rect 46293 44863 46351 44869
rect 46293 44860 46305 44863
rect 45879 44832 46305 44860
rect 45879 44829 45891 44832
rect 45833 44823 45891 44829
rect 46293 44829 46305 44832
rect 46339 44829 46351 44863
rect 46293 44823 46351 44829
rect 9582 44792 9588 44804
rect 9495 44764 9588 44792
rect 9582 44752 9588 44764
rect 9640 44792 9646 44804
rect 22830 44792 22836 44804
rect 9640 44764 22836 44792
rect 9640 44752 9646 44764
rect 22830 44752 22836 44764
rect 22888 44752 22894 44804
rect 46474 44792 46480 44804
rect 46435 44764 46480 44792
rect 46474 44752 46480 44764
rect 46532 44752 46538 44804
rect 38286 44684 38292 44736
rect 38344 44724 38350 44736
rect 47578 44724 47584 44736
rect 38344 44696 47584 44724
rect 38344 44684 38350 44696
rect 47578 44684 47584 44696
rect 47636 44684 47642 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 3050 44480 3056 44532
rect 3108 44520 3114 44532
rect 15562 44520 15568 44532
rect 3108 44492 15568 44520
rect 3108 44480 3114 44492
rect 15562 44480 15568 44492
rect 15620 44480 15626 44532
rect 46293 44523 46351 44529
rect 46293 44489 46305 44523
rect 46339 44520 46351 44523
rect 46474 44520 46480 44532
rect 46339 44492 46480 44520
rect 46339 44489 46351 44492
rect 46293 44483 46351 44489
rect 46474 44480 46480 44492
rect 46532 44480 46538 44532
rect 29914 44412 29920 44464
rect 29972 44452 29978 44464
rect 29972 44424 47624 44452
rect 29972 44412 29978 44424
rect 9125 44387 9183 44393
rect 9125 44353 9137 44387
rect 9171 44384 9183 44387
rect 9214 44384 9220 44396
rect 9171 44356 9220 44384
rect 9171 44353 9183 44356
rect 9125 44347 9183 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 38010 44344 38016 44396
rect 38068 44384 38074 44396
rect 47596 44393 47624 44424
rect 46201 44387 46259 44393
rect 46201 44384 46213 44387
rect 38068 44356 46213 44384
rect 38068 44344 38074 44356
rect 46201 44353 46213 44356
rect 46247 44353 46259 44387
rect 46201 44347 46259 44353
rect 47581 44387 47639 44393
rect 47581 44353 47593 44387
rect 47627 44384 47639 44387
rect 47854 44384 47860 44396
rect 47627 44356 47860 44384
rect 47627 44353 47639 44356
rect 47581 44347 47639 44353
rect 47854 44344 47860 44356
rect 47912 44344 47918 44396
rect 9030 44276 9036 44328
rect 9088 44316 9094 44328
rect 9401 44319 9459 44325
rect 9401 44316 9413 44319
rect 9088 44288 9413 44316
rect 9088 44276 9094 44288
rect 9401 44285 9413 44288
rect 9447 44316 9459 44319
rect 32766 44316 32772 44328
rect 9447 44288 32772 44316
rect 9447 44285 9459 44288
rect 9401 44279 9459 44285
rect 32766 44276 32772 44288
rect 32824 44276 32830 44328
rect 45370 44208 45376 44260
rect 45428 44248 45434 44260
rect 47673 44251 47731 44257
rect 47673 44248 47685 44251
rect 45428 44220 47685 44248
rect 45428 44208 45434 44220
rect 47673 44217 47685 44220
rect 47719 44217 47731 44251
rect 47673 44211 47731 44217
rect 45186 44140 45192 44192
rect 45244 44180 45250 44192
rect 47029 44183 47087 44189
rect 47029 44180 47041 44183
rect 45244 44152 47041 44180
rect 45244 44140 45250 44152
rect 47029 44149 47041 44152
rect 47075 44149 47087 44183
rect 47029 44143 47087 44149
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 48038 43840 48044 43852
rect 47999 43812 48044 43840
rect 48038 43800 48044 43812
rect 48096 43800 48102 43852
rect 2130 43732 2136 43784
rect 2188 43772 2194 43784
rect 2317 43775 2375 43781
rect 2317 43772 2329 43775
rect 2188 43744 2329 43772
rect 2188 43732 2194 43744
rect 2317 43741 2329 43744
rect 2363 43741 2375 43775
rect 2317 43735 2375 43741
rect 40034 43732 40040 43784
rect 40092 43772 40098 43784
rect 40405 43775 40463 43781
rect 40405 43772 40417 43775
rect 40092 43744 40417 43772
rect 40092 43732 40098 43744
rect 40405 43741 40417 43744
rect 40451 43741 40463 43775
rect 40405 43735 40463 43741
rect 46014 43732 46020 43784
rect 46072 43772 46078 43784
rect 46293 43775 46351 43781
rect 46293 43772 46305 43775
rect 46072 43744 46305 43772
rect 46072 43732 46078 43744
rect 46293 43741 46305 43744
rect 46339 43741 46351 43775
rect 46293 43735 46351 43741
rect 46477 43707 46535 43713
rect 46477 43673 46489 43707
rect 46523 43704 46535 43707
rect 46566 43704 46572 43716
rect 46523 43676 46572 43704
rect 46523 43673 46535 43676
rect 46477 43667 46535 43673
rect 46566 43664 46572 43676
rect 46624 43664 46630 43716
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 46566 43432 46572 43444
rect 46527 43404 46572 43432
rect 46566 43392 46572 43404
rect 46624 43392 46630 43444
rect 3970 43364 3976 43376
rect 3931 43336 3976 43364
rect 3970 43324 3976 43336
rect 4028 43324 4034 43376
rect 2130 43296 2136 43308
rect 2091 43268 2136 43296
rect 2130 43256 2136 43268
rect 2188 43256 2194 43308
rect 40034 43296 40040 43308
rect 39995 43268 40040 43296
rect 40034 43256 40040 43268
rect 40092 43256 40098 43308
rect 46014 43296 46020 43308
rect 45975 43268 46020 43296
rect 46014 43256 46020 43268
rect 46072 43256 46078 43308
rect 46474 43296 46480 43308
rect 46435 43268 46480 43296
rect 46474 43256 46480 43268
rect 46532 43256 46538 43308
rect 47578 43296 47584 43308
rect 47539 43268 47584 43296
rect 47578 43256 47584 43268
rect 47636 43256 47642 43308
rect 2317 43231 2375 43237
rect 2317 43197 2329 43231
rect 2363 43228 2375 43231
rect 3878 43228 3884 43240
rect 2363 43200 3884 43228
rect 2363 43197 2375 43200
rect 2317 43191 2375 43197
rect 3878 43188 3884 43200
rect 3936 43188 3942 43240
rect 40218 43228 40224 43240
rect 40179 43200 40224 43228
rect 40218 43188 40224 43200
rect 40276 43188 40282 43240
rect 41414 43228 41420 43240
rect 41375 43200 41420 43228
rect 41414 43188 41420 43200
rect 41472 43188 41478 43240
rect 47670 43092 47676 43104
rect 47631 43064 47676 43092
rect 47670 43052 47676 43064
rect 47728 43052 47734 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 3878 42752 3884 42764
rect 3839 42724 3884 42752
rect 3878 42712 3884 42724
rect 3936 42712 3942 42764
rect 26973 42755 27031 42761
rect 26973 42721 26985 42755
rect 27019 42752 27031 42755
rect 27985 42755 28043 42761
rect 27985 42752 27997 42755
rect 27019 42724 27997 42752
rect 27019 42721 27031 42724
rect 26973 42715 27031 42721
rect 27985 42721 27997 42724
rect 28031 42752 28043 42755
rect 30650 42752 30656 42764
rect 28031 42724 30656 42752
rect 28031 42721 28043 42724
rect 27985 42715 28043 42721
rect 30650 42712 30656 42724
rect 30708 42712 30714 42764
rect 46477 42755 46535 42761
rect 46477 42721 46489 42755
rect 46523 42752 46535 42755
rect 47670 42752 47676 42764
rect 46523 42724 47676 42752
rect 46523 42721 46535 42724
rect 46477 42715 46535 42721
rect 47670 42712 47676 42724
rect 47728 42712 47734 42764
rect 3789 42687 3847 42693
rect 3789 42653 3801 42687
rect 3835 42684 3847 42687
rect 6362 42684 6368 42696
rect 3835 42656 6368 42684
rect 3835 42653 3847 42656
rect 3789 42647 3847 42653
rect 6362 42644 6368 42656
rect 6420 42684 6426 42696
rect 9582 42684 9588 42696
rect 6420 42656 9588 42684
rect 6420 42644 6426 42656
rect 9582 42644 9588 42656
rect 9640 42644 9646 42696
rect 27157 42687 27215 42693
rect 27157 42653 27169 42687
rect 27203 42684 27215 42687
rect 27614 42684 27620 42696
rect 27203 42656 27620 42684
rect 27203 42653 27215 42656
rect 27157 42647 27215 42653
rect 27614 42644 27620 42656
rect 27672 42644 27678 42696
rect 28169 42687 28227 42693
rect 28169 42653 28181 42687
rect 28215 42653 28227 42687
rect 28169 42647 28227 42653
rect 33689 42687 33747 42693
rect 33689 42653 33701 42687
rect 33735 42684 33747 42687
rect 33778 42684 33784 42696
rect 33735 42656 33784 42684
rect 33735 42653 33747 42656
rect 33689 42647 33747 42653
rect 8938 42576 8944 42628
rect 8996 42616 9002 42628
rect 27709 42619 27767 42625
rect 27709 42616 27721 42619
rect 8996 42588 27721 42616
rect 8996 42576 9002 42588
rect 27709 42585 27721 42588
rect 27755 42616 27767 42619
rect 28184 42616 28212 42647
rect 33778 42644 33784 42656
rect 33836 42644 33842 42696
rect 45189 42687 45247 42693
rect 45189 42653 45201 42687
rect 45235 42684 45247 42687
rect 45738 42684 45744 42696
rect 45235 42656 45744 42684
rect 45235 42653 45247 42656
rect 45189 42647 45247 42653
rect 45738 42644 45744 42656
rect 45796 42644 45802 42696
rect 45833 42687 45891 42693
rect 45833 42653 45845 42687
rect 45879 42684 45891 42687
rect 46293 42687 46351 42693
rect 46293 42684 46305 42687
rect 45879 42656 46305 42684
rect 45879 42653 45891 42656
rect 45833 42647 45891 42653
rect 46293 42653 46305 42656
rect 46339 42653 46351 42687
rect 46293 42647 46351 42653
rect 48130 42616 48136 42628
rect 27755 42588 28212 42616
rect 48091 42588 48136 42616
rect 27755 42585 27767 42588
rect 27709 42579 27767 42585
rect 48130 42576 48136 42588
rect 48188 42576 48194 42628
rect 27154 42508 27160 42560
rect 27212 42548 27218 42560
rect 27341 42551 27399 42557
rect 27341 42548 27353 42551
rect 27212 42520 27353 42548
rect 27212 42508 27218 42520
rect 27341 42517 27353 42520
rect 27387 42517 27399 42551
rect 27341 42511 27399 42517
rect 28353 42551 28411 42557
rect 28353 42517 28365 42551
rect 28399 42548 28411 42551
rect 28534 42548 28540 42560
rect 28399 42520 28540 42548
rect 28399 42517 28411 42520
rect 28353 42511 28411 42517
rect 28534 42508 28540 42520
rect 28592 42508 28598 42560
rect 33502 42548 33508 42560
rect 33463 42520 33508 42548
rect 33502 42508 33508 42520
rect 33560 42508 33566 42560
rect 45005 42551 45063 42557
rect 45005 42517 45017 42551
rect 45051 42548 45063 42551
rect 45278 42548 45284 42560
rect 45051 42520 45284 42548
rect 45051 42517 45063 42520
rect 45005 42511 45063 42517
rect 45278 42508 45284 42520
rect 45336 42508 45342 42560
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 40218 42304 40224 42356
rect 40276 42344 40282 42356
rect 40313 42347 40371 42353
rect 40313 42344 40325 42347
rect 40276 42316 40325 42344
rect 40276 42304 40282 42316
rect 40313 42313 40325 42316
rect 40359 42313 40371 42347
rect 40313 42307 40371 42313
rect 33404 42279 33462 42285
rect 33404 42245 33416 42279
rect 33450 42276 33462 42279
rect 33502 42276 33508 42288
rect 33450 42248 33508 42276
rect 33450 42245 33462 42248
rect 33404 42239 33462 42245
rect 33502 42236 33508 42248
rect 33560 42236 33566 42288
rect 37645 42279 37703 42285
rect 37645 42276 37657 42279
rect 36648 42248 37657 42276
rect 27154 42208 27160 42220
rect 27115 42180 27160 42208
rect 27154 42168 27160 42180
rect 27212 42168 27218 42220
rect 28534 42208 28540 42220
rect 28495 42180 28540 42208
rect 28534 42168 28540 42180
rect 28592 42168 28598 42220
rect 31386 42208 31392 42220
rect 31347 42180 31392 42208
rect 31386 42168 31392 42180
rect 31444 42168 31450 42220
rect 32674 42208 32680 42220
rect 32635 42180 32680 42208
rect 32674 42168 32680 42180
rect 32732 42168 32738 42220
rect 36648 42217 36676 42248
rect 37645 42245 37657 42248
rect 37691 42245 37703 42279
rect 45370 42276 45376 42288
rect 45331 42248 45376 42276
rect 37645 42239 37703 42245
rect 45370 42236 45376 42248
rect 45428 42236 45434 42288
rect 35161 42211 35219 42217
rect 35161 42177 35173 42211
rect 35207 42177 35219 42211
rect 35161 42171 35219 42177
rect 35345 42211 35403 42217
rect 35345 42177 35357 42211
rect 35391 42208 35403 42211
rect 35989 42211 36047 42217
rect 35989 42208 36001 42211
rect 35391 42180 36001 42208
rect 35391 42177 35403 42180
rect 35345 42171 35403 42177
rect 35989 42177 36001 42180
rect 36035 42177 36047 42211
rect 35989 42171 36047 42177
rect 36633 42211 36691 42217
rect 36633 42177 36645 42211
rect 36679 42177 36691 42211
rect 36633 42171 36691 42177
rect 37461 42211 37519 42217
rect 37461 42177 37473 42211
rect 37507 42208 37519 42211
rect 38194 42208 38200 42220
rect 37507 42180 38200 42208
rect 37507 42177 37519 42180
rect 37461 42171 37519 42177
rect 33134 42140 33140 42152
rect 33095 42112 33140 42140
rect 33134 42100 33140 42112
rect 33192 42100 33198 42152
rect 34977 42143 35035 42149
rect 34977 42109 34989 42143
rect 35023 42109 35035 42143
rect 34977 42103 35035 42109
rect 26970 42004 26976 42016
rect 26931 41976 26976 42004
rect 26970 41964 26976 41976
rect 27028 41964 27034 42016
rect 28353 42007 28411 42013
rect 28353 41973 28365 42007
rect 28399 42004 28411 42007
rect 29638 42004 29644 42016
rect 28399 41976 29644 42004
rect 28399 41973 28411 41976
rect 28353 41967 28411 41973
rect 29638 41964 29644 41976
rect 29696 41964 29702 42016
rect 31202 42004 31208 42016
rect 31163 41976 31208 42004
rect 31202 41964 31208 41976
rect 31260 41964 31266 42016
rect 32490 42004 32496 42016
rect 32451 41976 32496 42004
rect 32490 41964 32496 41976
rect 32548 41964 32554 42016
rect 34514 42004 34520 42016
rect 34427 41976 34520 42004
rect 34514 41964 34520 41976
rect 34572 42004 34578 42016
rect 34992 42004 35020 42103
rect 35176 42072 35204 42171
rect 36722 42100 36728 42152
rect 36780 42140 36786 42152
rect 37277 42143 37335 42149
rect 37277 42140 37289 42143
rect 36780 42112 37289 42140
rect 36780 42100 36786 42112
rect 37277 42109 37289 42112
rect 37323 42109 37335 42143
rect 37277 42103 37335 42109
rect 37476 42072 37504 42171
rect 38194 42168 38200 42180
rect 38252 42168 38258 42220
rect 40221 42211 40279 42217
rect 40221 42177 40233 42211
rect 40267 42208 40279 42211
rect 41138 42208 41144 42220
rect 40267 42180 41144 42208
rect 40267 42177 40279 42180
rect 40221 42171 40279 42177
rect 41138 42168 41144 42180
rect 41196 42168 41202 42220
rect 41598 42208 41604 42220
rect 41559 42180 41604 42208
rect 41598 42168 41604 42180
rect 41656 42168 41662 42220
rect 41693 42211 41751 42217
rect 41693 42177 41705 42211
rect 41739 42177 41751 42211
rect 42518 42208 42524 42220
rect 42479 42180 42524 42208
rect 41693 42171 41751 42177
rect 41708 42140 41736 42171
rect 42518 42168 42524 42180
rect 42576 42168 42582 42220
rect 42613 42211 42671 42217
rect 42613 42177 42625 42211
rect 42659 42177 42671 42211
rect 42613 42171 42671 42177
rect 42797 42211 42855 42217
rect 42797 42177 42809 42211
rect 42843 42208 42855 42211
rect 43441 42211 43499 42217
rect 43441 42208 43453 42211
rect 42843 42180 43453 42208
rect 42843 42177 42855 42180
rect 42797 42171 42855 42177
rect 43441 42177 43453 42180
rect 43487 42177 43499 42211
rect 45186 42208 45192 42220
rect 45147 42180 45192 42208
rect 43441 42171 43499 42177
rect 42628 42140 42656 42171
rect 45186 42168 45192 42180
rect 45244 42168 45250 42220
rect 46842 42140 46848 42152
rect 40236 42112 42656 42140
rect 46803 42112 46848 42140
rect 40236 42084 40264 42112
rect 46842 42100 46848 42112
rect 46900 42100 46906 42152
rect 35176 42044 37504 42072
rect 40218 42032 40224 42084
rect 40276 42032 40282 42084
rect 35342 42004 35348 42016
rect 34572 41976 35348 42004
rect 34572 41964 34578 41976
rect 35342 41964 35348 41976
rect 35400 41964 35406 42016
rect 35802 42004 35808 42016
rect 35763 41976 35808 42004
rect 35802 41964 35808 41976
rect 35860 41964 35866 42016
rect 36446 42004 36452 42016
rect 36407 41976 36452 42004
rect 36446 41964 36452 41976
rect 36504 41964 36510 42016
rect 41874 42004 41880 42016
rect 41835 41976 41880 42004
rect 41874 41964 41880 41976
rect 41932 41964 41938 42016
rect 43254 42004 43260 42016
rect 43215 41976 43260 42004
rect 43254 41964 43260 41976
rect 43312 41964 43318 42016
rect 46290 41964 46296 42016
rect 46348 42004 46354 42016
rect 47765 42007 47823 42013
rect 47765 42004 47777 42007
rect 46348 41976 47777 42004
rect 46348 41964 46354 41976
rect 47765 41973 47777 41976
rect 47811 41973 47823 42007
rect 47765 41967 47823 41973
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 32674 41760 32680 41812
rect 32732 41800 32738 41812
rect 33597 41803 33655 41809
rect 33597 41800 33609 41803
rect 32732 41772 33609 41800
rect 32732 41760 32738 41772
rect 33597 41769 33609 41772
rect 33643 41769 33655 41803
rect 33597 41763 33655 41769
rect 36633 41803 36691 41809
rect 36633 41769 36645 41803
rect 36679 41800 36691 41803
rect 36722 41800 36728 41812
rect 36679 41772 36728 41800
rect 36679 41769 36691 41772
rect 36633 41763 36691 41769
rect 36722 41760 36728 41772
rect 36780 41760 36786 41812
rect 42518 41800 42524 41812
rect 42479 41772 42524 41800
rect 42518 41760 42524 41772
rect 42576 41760 42582 41812
rect 35253 41667 35311 41673
rect 35253 41664 35265 41667
rect 33152 41636 35265 41664
rect 33152 41608 33180 41636
rect 35253 41633 35265 41636
rect 35299 41633 35311 41667
rect 40218 41664 40224 41676
rect 35253 41627 35311 41633
rect 40052 41636 40224 41664
rect 26513 41599 26571 41605
rect 26513 41565 26525 41599
rect 26559 41596 26571 41599
rect 29546 41596 29552 41608
rect 26559 41568 29552 41596
rect 26559 41565 26571 41568
rect 26513 41559 26571 41565
rect 29546 41556 29552 41568
rect 29604 41556 29610 41608
rect 29638 41556 29644 41608
rect 29696 41596 29702 41608
rect 29805 41599 29863 41605
rect 29805 41596 29817 41599
rect 29696 41568 29817 41596
rect 29696 41556 29702 41568
rect 29805 41565 29817 41568
rect 29851 41565 29863 41599
rect 29805 41559 29863 41565
rect 31389 41599 31447 41605
rect 31389 41565 31401 41599
rect 31435 41596 31447 41599
rect 33134 41596 33140 41608
rect 31435 41568 33140 41596
rect 31435 41565 31447 41568
rect 31389 41559 31447 41565
rect 33134 41556 33140 41568
rect 33192 41556 33198 41608
rect 33321 41599 33379 41605
rect 33321 41565 33333 41599
rect 33367 41565 33379 41599
rect 33321 41559 33379 41565
rect 33413 41599 33471 41605
rect 33413 41565 33425 41599
rect 33459 41596 33471 41599
rect 33594 41596 33600 41608
rect 33459 41568 33600 41596
rect 33459 41565 33471 41568
rect 33413 41559 33471 41565
rect 26780 41531 26838 41537
rect 26780 41497 26792 41531
rect 26826 41528 26838 41531
rect 26970 41528 26976 41540
rect 26826 41500 26976 41528
rect 26826 41497 26838 41500
rect 26780 41491 26838 41497
rect 26970 41488 26976 41500
rect 27028 41488 27034 41540
rect 31202 41488 31208 41540
rect 31260 41528 31266 41540
rect 31634 41531 31692 41537
rect 31634 41528 31646 41531
rect 31260 41500 31646 41528
rect 31260 41488 31266 41500
rect 31634 41497 31646 41500
rect 31680 41497 31692 41531
rect 33336 41528 33364 41559
rect 33594 41556 33600 41568
rect 33652 41556 33658 41608
rect 35520 41599 35578 41605
rect 35520 41565 35532 41599
rect 35566 41596 35578 41599
rect 35802 41596 35808 41608
rect 35566 41568 35808 41596
rect 35566 41565 35578 41568
rect 35520 41559 35578 41565
rect 35802 41556 35808 41568
rect 35860 41556 35866 41608
rect 37093 41599 37151 41605
rect 37093 41565 37105 41599
rect 37139 41596 37151 41599
rect 37642 41596 37648 41608
rect 37139 41568 37648 41596
rect 37139 41565 37151 41568
rect 37093 41559 37151 41565
rect 37642 41556 37648 41568
rect 37700 41556 37706 41608
rect 39301 41599 39359 41605
rect 39301 41565 39313 41599
rect 39347 41565 39359 41599
rect 39301 41559 39359 41565
rect 34606 41528 34612 41540
rect 31634 41491 31692 41497
rect 32784 41500 34612 41528
rect 27890 41460 27896 41472
rect 27851 41432 27896 41460
rect 27890 41420 27896 41432
rect 27948 41420 27954 41472
rect 30926 41460 30932 41472
rect 30887 41432 30932 41460
rect 30926 41420 30932 41432
rect 30984 41420 30990 41472
rect 32784 41469 32812 41500
rect 34606 41488 34612 41500
rect 34664 41488 34670 41540
rect 36446 41488 36452 41540
rect 36504 41528 36510 41540
rect 37338 41531 37396 41537
rect 37338 41528 37350 41531
rect 36504 41500 37350 41528
rect 36504 41488 36510 41500
rect 37338 41497 37350 41500
rect 37384 41497 37396 41531
rect 39316 41528 39344 41559
rect 39390 41556 39396 41608
rect 39448 41596 39454 41608
rect 40052 41605 40080 41636
rect 40218 41624 40224 41636
rect 40276 41624 40282 41676
rect 46290 41664 46296 41676
rect 46251 41636 46296 41664
rect 46290 41624 46296 41636
rect 46348 41624 46354 41676
rect 39853 41599 39911 41605
rect 39853 41596 39865 41599
rect 39448 41568 39865 41596
rect 39448 41556 39454 41568
rect 39853 41565 39865 41568
rect 39899 41565 39911 41599
rect 39853 41559 39911 41565
rect 40037 41599 40095 41605
rect 40037 41565 40049 41599
rect 40083 41565 40095 41599
rect 40037 41559 40095 41565
rect 40126 41556 40132 41608
rect 40184 41596 40190 41608
rect 41141 41599 41199 41605
rect 41141 41596 41153 41599
rect 40184 41568 41153 41596
rect 40184 41556 40190 41568
rect 41141 41565 41153 41568
rect 41187 41565 41199 41599
rect 41141 41559 41199 41565
rect 42981 41599 43039 41605
rect 42981 41565 42993 41599
rect 43027 41596 43039 41599
rect 43990 41596 43996 41608
rect 43027 41568 43996 41596
rect 43027 41565 43039 41568
rect 42981 41559 43039 41565
rect 43990 41556 43996 41568
rect 44048 41556 44054 41608
rect 45094 41596 45100 41608
rect 45055 41568 45100 41596
rect 45094 41556 45100 41568
rect 45152 41556 45158 41608
rect 45278 41596 45284 41608
rect 45239 41568 45284 41596
rect 45278 41556 45284 41568
rect 45336 41556 45342 41608
rect 40221 41531 40279 41537
rect 40221 41528 40233 41531
rect 39316 41500 40233 41528
rect 37338 41491 37396 41497
rect 40221 41497 40233 41500
rect 40267 41497 40279 41531
rect 40221 41491 40279 41497
rect 41408 41531 41466 41537
rect 41408 41497 41420 41531
rect 41454 41528 41466 41531
rect 41690 41528 41696 41540
rect 41454 41500 41696 41528
rect 41454 41497 41466 41500
rect 41408 41491 41466 41497
rect 41690 41488 41696 41500
rect 41748 41488 41754 41540
rect 43254 41537 43260 41540
rect 43248 41528 43260 41537
rect 43215 41500 43260 41528
rect 43248 41491 43260 41500
rect 43254 41488 43260 41491
rect 43312 41488 43318 41540
rect 46477 41531 46535 41537
rect 46477 41497 46489 41531
rect 46523 41528 46535 41531
rect 46934 41528 46940 41540
rect 46523 41500 46940 41528
rect 46523 41497 46535 41500
rect 46477 41491 46535 41497
rect 46934 41488 46940 41500
rect 46992 41488 46998 41540
rect 48133 41531 48191 41537
rect 48133 41497 48145 41531
rect 48179 41528 48191 41531
rect 48222 41528 48228 41540
rect 48179 41500 48228 41528
rect 48179 41497 48191 41500
rect 48133 41491 48191 41497
rect 48222 41488 48228 41500
rect 48280 41488 48286 41540
rect 32769 41463 32827 41469
rect 32769 41429 32781 41463
rect 32815 41429 32827 41463
rect 32769 41423 32827 41429
rect 38102 41420 38108 41472
rect 38160 41460 38166 41472
rect 38473 41463 38531 41469
rect 38473 41460 38485 41463
rect 38160 41432 38485 41460
rect 38160 41420 38166 41432
rect 38473 41429 38485 41432
rect 38519 41429 38531 41463
rect 38473 41423 38531 41429
rect 39117 41463 39175 41469
rect 39117 41429 39129 41463
rect 39163 41460 39175 41463
rect 40034 41460 40040 41472
rect 39163 41432 40040 41460
rect 39163 41429 39175 41432
rect 39117 41423 39175 41429
rect 40034 41420 40040 41432
rect 40092 41420 40098 41472
rect 43806 41420 43812 41472
rect 43864 41460 43870 41472
rect 44361 41463 44419 41469
rect 44361 41460 44373 41463
rect 43864 41432 44373 41460
rect 43864 41420 43870 41432
rect 44361 41429 44373 41432
rect 44407 41429 44419 41463
rect 44361 41423 44419 41429
rect 45465 41463 45523 41469
rect 45465 41429 45477 41463
rect 45511 41460 45523 41463
rect 46014 41460 46020 41472
rect 45511 41432 46020 41460
rect 45511 41429 45523 41432
rect 45465 41423 45523 41429
rect 46014 41420 46020 41432
rect 46072 41420 46078 41472
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 31205 41259 31263 41265
rect 31205 41225 31217 41259
rect 31251 41256 31263 41259
rect 31386 41256 31392 41268
rect 31251 41228 31392 41256
rect 31251 41225 31263 41228
rect 31205 41219 31263 41225
rect 31386 41216 31392 41228
rect 31444 41216 31450 41268
rect 34422 41256 34428 41268
rect 32876 41228 34428 41256
rect 9033 41191 9091 41197
rect 9033 41157 9045 41191
rect 9079 41188 9091 41191
rect 17037 41191 17095 41197
rect 17037 41188 17049 41191
rect 9079 41160 17049 41188
rect 9079 41157 9091 41160
rect 9033 41151 9091 41157
rect 17037 41157 17049 41160
rect 17083 41157 17095 41191
rect 17037 41151 17095 41157
rect 32490 41148 32496 41200
rect 32548 41188 32554 41200
rect 32646 41191 32704 41197
rect 32646 41188 32658 41191
rect 32548 41160 32658 41188
rect 32548 41148 32554 41160
rect 32646 41157 32658 41160
rect 32692 41157 32704 41191
rect 32646 41151 32704 41157
rect 16942 41120 16948 41132
rect 16903 41092 16948 41120
rect 16942 41080 16948 41092
rect 17000 41080 17006 41132
rect 25501 41123 25559 41129
rect 25501 41089 25513 41123
rect 25547 41120 25559 41123
rect 26145 41123 26203 41129
rect 25547 41092 26096 41120
rect 25547 41089 25559 41092
rect 25501 41083 25559 41089
rect 8846 41052 8852 41064
rect 8807 41024 8852 41052
rect 8846 41012 8852 41024
rect 8904 41012 8910 41064
rect 9309 41055 9367 41061
rect 9309 41021 9321 41055
rect 9355 41021 9367 41055
rect 25958 41052 25964 41064
rect 25919 41024 25964 41052
rect 9309 41015 9367 41021
rect 3418 40944 3424 40996
rect 3476 40984 3482 40996
rect 9324 40984 9352 41015
rect 25958 41012 25964 41024
rect 26016 41012 26022 41064
rect 26068 41052 26096 41092
rect 26145 41089 26157 41123
rect 26191 41120 26203 41123
rect 27062 41120 27068 41132
rect 26191 41092 27068 41120
rect 26191 41089 26203 41092
rect 26145 41083 26203 41089
rect 27062 41080 27068 41092
rect 27120 41080 27126 41132
rect 28994 41080 29000 41132
rect 29052 41120 29058 41132
rect 29549 41123 29607 41129
rect 29549 41120 29561 41123
rect 29052 41092 29561 41120
rect 29052 41080 29058 41092
rect 29549 41089 29561 41092
rect 29595 41089 29607 41123
rect 29549 41083 29607 41089
rect 30006 41080 30012 41132
rect 30064 41120 30070 41132
rect 31021 41123 31079 41129
rect 31021 41120 31033 41123
rect 30064 41092 31033 41120
rect 30064 41080 30070 41092
rect 31021 41089 31033 41092
rect 31067 41089 31079 41123
rect 32876 41120 32904 41228
rect 34422 41216 34428 41228
rect 34480 41216 34486 41268
rect 39390 41256 39396 41268
rect 37384 41228 39396 41256
rect 37384 41200 37412 41228
rect 39390 41216 39396 41228
rect 39448 41216 39454 41268
rect 40034 41216 40040 41268
rect 40092 41256 40098 41268
rect 41690 41256 41696 41268
rect 40092 41228 40172 41256
rect 41651 41228 41696 41256
rect 40092 41216 40098 41228
rect 34514 41148 34520 41200
rect 34572 41188 34578 41200
rect 34572 41160 34617 41188
rect 34572 41148 34578 41160
rect 34698 41148 34704 41200
rect 34756 41188 34762 41200
rect 36265 41191 36323 41197
rect 34756 41160 35572 41188
rect 34756 41148 34762 41160
rect 31021 41083 31079 41089
rect 32324 41092 32904 41120
rect 34609 41123 34667 41129
rect 26602 41052 26608 41064
rect 26068 41024 26608 41052
rect 26602 41012 26608 41024
rect 26660 41012 26666 41064
rect 30837 41055 30895 41061
rect 30837 41021 30849 41055
rect 30883 41052 30895 41055
rect 30926 41052 30932 41064
rect 30883 41024 30932 41052
rect 30883 41021 30895 41024
rect 30837 41015 30895 41021
rect 30926 41012 30932 41024
rect 30984 41052 30990 41064
rect 32324 41052 32352 41092
rect 34609 41089 34621 41123
rect 34655 41118 34667 41123
rect 34790 41120 34796 41132
rect 34703 41118 34796 41120
rect 34655 41092 34796 41118
rect 34655 41090 34744 41092
rect 34655 41089 34667 41090
rect 34609 41083 34667 41089
rect 34790 41080 34796 41092
rect 34848 41120 34854 41132
rect 35544 41129 35572 41160
rect 36265 41157 36277 41191
rect 36311 41188 36323 41191
rect 37366 41188 37372 41200
rect 36311 41160 37372 41188
rect 36311 41157 36323 41160
rect 36265 41151 36323 41157
rect 37366 41148 37372 41160
rect 37424 41148 37430 41200
rect 37642 41148 37648 41200
rect 37700 41188 37706 41200
rect 40144 41197 40172 41228
rect 41690 41216 41696 41228
rect 41748 41216 41754 41268
rect 42705 41259 42763 41265
rect 42705 41225 42717 41259
rect 42751 41256 42763 41259
rect 42978 41256 42984 41268
rect 42751 41228 42984 41256
rect 42751 41225 42763 41228
rect 42705 41219 42763 41225
rect 42978 41216 42984 41228
rect 43036 41256 43042 41268
rect 45373 41259 45431 41265
rect 45373 41256 45385 41259
rect 43036 41228 45385 41256
rect 43036 41216 43042 41228
rect 45373 41225 45385 41228
rect 45419 41225 45431 41259
rect 46934 41256 46940 41268
rect 46895 41228 46940 41256
rect 45373 41219 45431 41225
rect 46934 41216 46940 41228
rect 46992 41216 46998 41268
rect 40120 41191 40178 41197
rect 37700 41160 39896 41188
rect 37700 41148 37706 41160
rect 35253 41123 35311 41129
rect 35253 41120 35265 41123
rect 34848 41092 35265 41120
rect 34848 41080 34854 41092
rect 35253 41089 35265 41092
rect 35299 41089 35311 41123
rect 35253 41083 35311 41089
rect 35529 41123 35587 41129
rect 35529 41089 35541 41123
rect 35575 41089 35587 41123
rect 35529 41083 35587 41089
rect 36541 41123 36599 41129
rect 36541 41089 36553 41123
rect 36587 41120 36599 41123
rect 36998 41120 37004 41132
rect 36587 41092 37004 41120
rect 36587 41089 36599 41092
rect 36541 41083 36599 41089
rect 36998 41080 37004 41092
rect 37056 41080 37062 41132
rect 37550 41120 37556 41132
rect 37511 41092 37556 41120
rect 37550 41080 37556 41092
rect 37608 41080 37614 41132
rect 38028 41129 38056 41160
rect 38013 41123 38071 41129
rect 38013 41089 38025 41123
rect 38059 41089 38071 41123
rect 38269 41123 38327 41129
rect 38269 41120 38281 41123
rect 38013 41083 38071 41089
rect 38120 41092 38281 41120
rect 30984 41024 32352 41052
rect 32401 41055 32459 41061
rect 30984 41012 30990 41024
rect 32401 41021 32413 41055
rect 32447 41021 32459 41055
rect 35342 41052 35348 41064
rect 35303 41024 35348 41052
rect 32401 41015 32459 41021
rect 3476 40956 9352 40984
rect 3476 40944 3482 40956
rect 24578 40944 24584 40996
rect 24636 40984 24642 40996
rect 26329 40987 26387 40993
rect 26329 40984 26341 40987
rect 24636 40956 26341 40984
rect 24636 40944 24642 40956
rect 26329 40953 26341 40956
rect 26375 40953 26387 40987
rect 26329 40947 26387 40953
rect 25314 40916 25320 40928
rect 25275 40888 25320 40916
rect 25314 40876 25320 40888
rect 25372 40876 25378 40928
rect 29362 40916 29368 40928
rect 29323 40888 29368 40916
rect 29362 40876 29368 40888
rect 29420 40876 29426 40928
rect 32416 40916 32444 41015
rect 35342 41012 35348 41024
rect 35400 41012 35406 41064
rect 36449 41055 36507 41061
rect 36449 41021 36461 41055
rect 36495 41052 36507 41055
rect 38120 41052 38148 41092
rect 38269 41089 38281 41092
rect 38315 41089 38327 41123
rect 38269 41083 38327 41089
rect 39868 41061 39896 41160
rect 40120 41157 40132 41191
rect 40166 41157 40178 41191
rect 40120 41151 40178 41157
rect 42429 41191 42487 41197
rect 42429 41157 42441 41191
rect 42475 41188 42487 41191
rect 42518 41188 42524 41200
rect 42475 41160 42524 41188
rect 42475 41157 42487 41160
rect 42429 41151 42487 41157
rect 42518 41148 42524 41160
rect 42576 41148 42582 41200
rect 41874 41120 41880 41132
rect 41835 41092 41880 41120
rect 41874 41080 41880 41092
rect 41932 41080 41938 41132
rect 42613 41123 42671 41129
rect 42613 41089 42625 41123
rect 42659 41089 42671 41123
rect 42613 41083 42671 41089
rect 42797 41123 42855 41129
rect 42797 41089 42809 41123
rect 42843 41120 42855 41123
rect 43806 41120 43812 41132
rect 42843 41092 43812 41120
rect 42843 41089 42855 41092
rect 42797 41083 42855 41089
rect 36495 41024 37320 41052
rect 36495 41021 36507 41024
rect 36449 41015 36507 41021
rect 33781 40987 33839 40993
rect 33781 40953 33793 40987
rect 33827 40984 33839 40987
rect 33870 40984 33876 40996
rect 33827 40956 33876 40984
rect 33827 40953 33839 40956
rect 33781 40947 33839 40953
rect 33870 40944 33876 40956
rect 33928 40944 33934 40996
rect 34241 40987 34299 40993
rect 34241 40953 34253 40987
rect 34287 40953 34299 40987
rect 34241 40947 34299 40953
rect 33134 40916 33140 40928
rect 32416 40888 33140 40916
rect 33134 40876 33140 40888
rect 33192 40916 33198 40928
rect 33686 40916 33692 40928
rect 33192 40888 33692 40916
rect 33192 40876 33198 40888
rect 33686 40876 33692 40888
rect 33744 40876 33750 40928
rect 34256 40916 34284 40947
rect 34422 40944 34428 40996
rect 34480 40984 34486 40996
rect 34480 40956 35296 40984
rect 34480 40944 34486 40956
rect 34606 40916 34612 40928
rect 34256 40888 34612 40916
rect 34606 40876 34612 40888
rect 34664 40876 34670 40928
rect 34790 40916 34796 40928
rect 34751 40888 34796 40916
rect 34790 40876 34796 40888
rect 34848 40876 34854 40928
rect 35268 40925 35296 40956
rect 35253 40919 35311 40925
rect 35253 40885 35265 40919
rect 35299 40885 35311 40919
rect 35710 40916 35716 40928
rect 35671 40888 35716 40916
rect 35253 40879 35311 40885
rect 35710 40876 35716 40888
rect 35768 40876 35774 40928
rect 36538 40916 36544 40928
rect 36499 40888 36544 40916
rect 36538 40876 36544 40888
rect 36596 40876 36602 40928
rect 36722 40916 36728 40928
rect 36683 40888 36728 40916
rect 36722 40876 36728 40888
rect 36780 40876 36786 40928
rect 37292 40916 37320 41024
rect 37384 41024 38148 41052
rect 39853 41055 39911 41061
rect 37384 40993 37412 41024
rect 39853 41021 39865 41055
rect 39899 41021 39911 41055
rect 39853 41015 39911 41021
rect 37369 40987 37427 40993
rect 37369 40953 37381 40987
rect 37415 40953 37427 40987
rect 37369 40947 37427 40953
rect 37458 40916 37464 40928
rect 37292 40888 37464 40916
rect 37458 40876 37464 40888
rect 37516 40876 37522 40928
rect 39868 40916 39896 41015
rect 41598 41012 41604 41064
rect 41656 41052 41662 41064
rect 42628 41052 42656 41083
rect 43806 41080 43812 41092
rect 43864 41080 43870 41132
rect 43990 41120 43996 41132
rect 43951 41092 43996 41120
rect 43990 41080 43996 41092
rect 44048 41080 44054 41132
rect 44082 41080 44088 41132
rect 44140 41120 44146 41132
rect 44249 41123 44307 41129
rect 44249 41120 44261 41123
rect 44140 41092 44261 41120
rect 44140 41080 44146 41092
rect 44249 41089 44261 41092
rect 44295 41089 44307 41123
rect 46014 41120 46020 41132
rect 45975 41092 46020 41120
rect 44249 41083 44307 41089
rect 46014 41080 46020 41092
rect 46072 41080 46078 41132
rect 46658 41080 46664 41132
rect 46716 41120 46722 41132
rect 46845 41123 46903 41129
rect 46845 41120 46857 41123
rect 46716 41092 46857 41120
rect 46716 41080 46722 41092
rect 46845 41089 46857 41092
rect 46891 41089 46903 41123
rect 46845 41083 46903 41089
rect 41656 41024 42656 41052
rect 41656 41012 41662 41024
rect 40126 40916 40132 40928
rect 39868 40888 40132 40916
rect 40126 40876 40132 40888
rect 40184 40876 40190 40928
rect 41230 40916 41236 40928
rect 41191 40888 41236 40916
rect 41230 40876 41236 40888
rect 41288 40876 41294 40928
rect 42794 40876 42800 40928
rect 42852 40916 42858 40928
rect 42981 40919 43039 40925
rect 42981 40916 42993 40919
rect 42852 40888 42993 40916
rect 42852 40876 42858 40888
rect 42981 40885 42993 40888
rect 43027 40885 43039 40919
rect 45830 40916 45836 40928
rect 45791 40888 45836 40916
rect 42981 40879 43039 40885
rect 45830 40876 45836 40888
rect 45888 40876 45894 40928
rect 46290 40876 46296 40928
rect 46348 40916 46354 40928
rect 47765 40919 47823 40925
rect 47765 40916 47777 40919
rect 46348 40888 47777 40916
rect 46348 40876 46354 40888
rect 47765 40885 47777 40888
rect 47811 40885 47823 40919
rect 47765 40879 47823 40885
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 8846 40672 8852 40724
rect 8904 40712 8910 40724
rect 9125 40715 9183 40721
rect 9125 40712 9137 40715
rect 8904 40684 9137 40712
rect 8904 40672 8910 40684
rect 9125 40681 9137 40684
rect 9171 40681 9183 40715
rect 9125 40675 9183 40681
rect 25958 40672 25964 40724
rect 26016 40712 26022 40724
rect 27890 40712 27896 40724
rect 26016 40684 27896 40712
rect 26016 40672 26022 40684
rect 27890 40672 27896 40684
rect 27948 40672 27954 40724
rect 28994 40712 29000 40724
rect 28955 40684 29000 40712
rect 28994 40672 29000 40684
rect 29052 40672 29058 40724
rect 32582 40712 32588 40724
rect 29564 40684 32588 40712
rect 27246 40604 27252 40656
rect 27304 40644 27310 40656
rect 29564 40644 29592 40684
rect 32582 40672 32588 40684
rect 32640 40672 32646 40724
rect 33778 40712 33784 40724
rect 33739 40684 33784 40712
rect 33778 40672 33784 40684
rect 33836 40672 33842 40724
rect 37550 40672 37556 40724
rect 37608 40712 37614 40724
rect 38381 40715 38439 40721
rect 38381 40712 38393 40715
rect 37608 40684 38393 40712
rect 37608 40672 37614 40684
rect 38381 40681 38393 40684
rect 38427 40681 38439 40715
rect 38381 40675 38439 40681
rect 38841 40715 38899 40721
rect 38841 40681 38853 40715
rect 38887 40712 38899 40715
rect 40218 40712 40224 40724
rect 38887 40684 40224 40712
rect 38887 40681 38899 40684
rect 38841 40675 38899 40681
rect 40218 40672 40224 40684
rect 40276 40712 40282 40724
rect 41598 40712 41604 40724
rect 40276 40684 41414 40712
rect 41559 40684 41604 40712
rect 40276 40672 40282 40684
rect 27304 40616 29592 40644
rect 27304 40604 27310 40616
rect 37642 40604 37648 40656
rect 37700 40644 37706 40656
rect 41386 40644 41414 40684
rect 41598 40672 41604 40684
rect 41656 40712 41662 40724
rect 42061 40715 42119 40721
rect 42061 40712 42073 40715
rect 41656 40684 42073 40712
rect 41656 40672 41662 40684
rect 42061 40681 42073 40684
rect 42107 40681 42119 40715
rect 42061 40675 42119 40681
rect 37700 40616 39068 40644
rect 41386 40616 43208 40644
rect 37700 40604 37706 40616
rect 2682 40536 2688 40588
rect 2740 40576 2746 40588
rect 22741 40579 22799 40585
rect 22741 40576 22753 40579
rect 2740 40548 22753 40576
rect 2740 40536 2746 40548
rect 22741 40545 22753 40548
rect 22787 40576 22799 40579
rect 28629 40579 28687 40585
rect 28629 40576 28641 40579
rect 22787 40548 23336 40576
rect 22787 40545 22799 40548
rect 22741 40539 22799 40545
rect 23308 40517 23336 40548
rect 27908 40548 28641 40576
rect 27908 40520 27936 40548
rect 28629 40545 28641 40548
rect 28675 40545 28687 40579
rect 29546 40576 29552 40588
rect 29507 40548 29552 40576
rect 28629 40539 28687 40545
rect 29546 40536 29552 40548
rect 29604 40536 29610 40588
rect 36722 40576 36728 40588
rect 34992 40548 36728 40576
rect 23201 40511 23259 40517
rect 23201 40477 23213 40511
rect 23247 40477 23259 40511
rect 23201 40471 23259 40477
rect 23293 40511 23351 40517
rect 23293 40477 23305 40511
rect 23339 40477 23351 40511
rect 24578 40508 24584 40520
rect 24539 40480 24584 40508
rect 23293 40471 23351 40477
rect 23216 40440 23244 40471
rect 24578 40468 24584 40480
rect 24636 40468 24642 40520
rect 24854 40468 24860 40520
rect 24912 40508 24918 40520
rect 25314 40517 25320 40520
rect 25041 40511 25099 40517
rect 25041 40508 25053 40511
rect 24912 40480 25053 40508
rect 24912 40468 24918 40480
rect 25041 40477 25053 40480
rect 25087 40477 25099 40511
rect 25308 40508 25320 40517
rect 25275 40480 25320 40508
rect 25041 40471 25099 40477
rect 25308 40471 25320 40480
rect 25314 40468 25320 40471
rect 25372 40468 25378 40520
rect 26973 40511 27031 40517
rect 26973 40477 26985 40511
rect 27019 40477 27031 40511
rect 26973 40471 27031 40477
rect 23842 40440 23848 40452
rect 23216 40412 23848 40440
rect 23842 40400 23848 40412
rect 23900 40400 23906 40452
rect 26988 40440 27016 40471
rect 27062 40468 27068 40520
rect 27120 40508 27126 40520
rect 27890 40508 27896 40520
rect 27120 40480 27165 40508
rect 27851 40480 27896 40508
rect 27120 40468 27126 40480
rect 27890 40468 27896 40480
rect 27948 40468 27954 40520
rect 27982 40468 27988 40520
rect 28040 40508 28046 40520
rect 28813 40511 28871 40517
rect 28040 40480 28085 40508
rect 28040 40468 28046 40480
rect 28813 40477 28825 40511
rect 28859 40508 28871 40511
rect 28859 40480 29316 40508
rect 28859 40477 28871 40480
rect 28813 40471 28871 40477
rect 27706 40440 27712 40452
rect 26436 40412 27712 40440
rect 23474 40372 23480 40384
rect 23435 40344 23480 40372
rect 23474 40332 23480 40344
rect 23532 40332 23538 40384
rect 24394 40372 24400 40384
rect 24355 40344 24400 40372
rect 24394 40332 24400 40344
rect 24452 40332 24458 40384
rect 26436 40381 26464 40412
rect 27706 40400 27712 40412
rect 27764 40400 27770 40452
rect 29178 40440 29184 40452
rect 28092 40412 29184 40440
rect 26421 40375 26479 40381
rect 26421 40341 26433 40375
rect 26467 40341 26479 40375
rect 26421 40335 26479 40341
rect 27249 40375 27307 40381
rect 27249 40341 27261 40375
rect 27295 40372 27307 40375
rect 28092 40372 28120 40412
rect 29178 40400 29184 40412
rect 29236 40400 29242 40452
rect 29288 40440 29316 40480
rect 29362 40468 29368 40520
rect 29420 40508 29426 40520
rect 29805 40511 29863 40517
rect 29805 40508 29817 40511
rect 29420 40480 29817 40508
rect 29420 40468 29426 40480
rect 29805 40477 29817 40480
rect 29851 40477 29863 40511
rect 29805 40471 29863 40477
rect 33505 40511 33563 40517
rect 33505 40477 33517 40511
rect 33551 40477 33563 40511
rect 33505 40471 33563 40477
rect 30006 40440 30012 40452
rect 29288 40412 30012 40440
rect 30006 40400 30012 40412
rect 30064 40400 30070 40452
rect 33520 40440 33548 40471
rect 33594 40468 33600 40520
rect 33652 40508 33658 40520
rect 34992 40517 35020 40548
rect 36722 40536 36728 40548
rect 36780 40536 36786 40588
rect 34977 40511 35035 40517
rect 33652 40480 34928 40508
rect 33652 40468 33658 40480
rect 33870 40440 33876 40452
rect 33520 40412 33876 40440
rect 33870 40400 33876 40412
rect 33928 40400 33934 40452
rect 34900 40440 34928 40480
rect 34977 40477 34989 40511
rect 35023 40477 35035 40511
rect 34977 40471 35035 40477
rect 35161 40511 35219 40517
rect 35161 40477 35173 40511
rect 35207 40508 35219 40511
rect 35710 40508 35716 40520
rect 35207 40480 35716 40508
rect 35207 40477 35219 40480
rect 35161 40471 35219 40477
rect 35710 40468 35716 40480
rect 35768 40468 35774 40520
rect 36541 40511 36599 40517
rect 36541 40477 36553 40511
rect 36587 40508 36599 40511
rect 36630 40508 36636 40520
rect 36587 40480 36636 40508
rect 36587 40477 36599 40480
rect 36541 40471 36599 40477
rect 36630 40468 36636 40480
rect 36688 40468 36694 40520
rect 36998 40508 37004 40520
rect 36911 40480 37004 40508
rect 36998 40468 37004 40480
rect 37056 40508 37062 40520
rect 37292 40508 37381 40510
rect 38102 40508 38108 40520
rect 37056 40482 38108 40508
rect 37056 40480 37320 40482
rect 37353 40480 38108 40482
rect 37056 40468 37062 40480
rect 38102 40468 38108 40480
rect 38160 40468 38166 40520
rect 38194 40468 38200 40520
rect 38252 40508 38258 40520
rect 39040 40517 39068 40616
rect 42245 40579 42303 40585
rect 42245 40545 42257 40579
rect 42291 40576 42303 40579
rect 42978 40576 42984 40588
rect 42291 40548 42984 40576
rect 42291 40545 42303 40548
rect 42245 40539 42303 40545
rect 42978 40536 42984 40548
rect 43036 40536 43042 40588
rect 43180 40576 43208 40616
rect 46290 40576 46296 40588
rect 43180 40548 44036 40576
rect 46251 40548 46296 40576
rect 39025 40511 39083 40517
rect 38252 40480 38297 40508
rect 38252 40468 38258 40480
rect 39025 40477 39037 40511
rect 39071 40477 39083 40511
rect 40218 40508 40224 40520
rect 40179 40480 40224 40508
rect 39025 40471 39083 40477
rect 40218 40468 40224 40480
rect 40276 40468 40282 40520
rect 42337 40511 42395 40517
rect 42337 40477 42349 40511
rect 42383 40508 42395 40511
rect 42518 40508 42524 40520
rect 42383 40480 42524 40508
rect 42383 40477 42395 40480
rect 42337 40471 42395 40477
rect 42518 40468 42524 40480
rect 42576 40468 42582 40520
rect 43180 40517 43208 40548
rect 43165 40511 43223 40517
rect 43165 40477 43177 40511
rect 43211 40477 43223 40511
rect 43806 40508 43812 40520
rect 43767 40480 43812 40508
rect 43165 40471 43223 40477
rect 43806 40468 43812 40480
rect 43864 40468 43870 40520
rect 44008 40517 44036 40548
rect 46290 40536 46296 40548
rect 46348 40536 46354 40588
rect 43993 40511 44051 40517
rect 43993 40477 44005 40511
rect 44039 40477 44051 40511
rect 43993 40471 44051 40477
rect 34900 40412 36400 40440
rect 36372 40384 36400 40412
rect 37366 40400 37372 40452
rect 37424 40440 37430 40452
rect 37550 40440 37556 40452
rect 37424 40412 37469 40440
rect 37511 40412 37556 40440
rect 37424 40400 37430 40412
rect 37550 40400 37556 40412
rect 37608 40400 37614 40452
rect 40488 40443 40546 40449
rect 40488 40409 40500 40443
rect 40534 40440 40546 40443
rect 40678 40440 40684 40452
rect 40534 40412 40684 40440
rect 40534 40409 40546 40412
rect 40488 40403 40546 40409
rect 40678 40400 40684 40412
rect 40736 40400 40742 40452
rect 42061 40443 42119 40449
rect 42061 40409 42073 40443
rect 42107 40440 42119 40443
rect 43824 40440 43852 40468
rect 42107 40412 43852 40440
rect 46477 40443 46535 40449
rect 42107 40409 42119 40412
rect 42061 40403 42119 40409
rect 46477 40409 46489 40443
rect 46523 40440 46535 40443
rect 46934 40440 46940 40452
rect 46523 40412 46940 40440
rect 46523 40409 46535 40412
rect 46477 40403 46535 40409
rect 46934 40400 46940 40412
rect 46992 40400 46998 40452
rect 48130 40440 48136 40452
rect 48091 40412 48136 40440
rect 48130 40400 48136 40412
rect 48188 40400 48194 40452
rect 27295 40344 28120 40372
rect 27295 40341 27307 40344
rect 27249 40335 27307 40341
rect 28166 40332 28172 40384
rect 28224 40372 28230 40384
rect 28224 40344 28269 40372
rect 28224 40332 28230 40344
rect 30742 40332 30748 40384
rect 30800 40372 30806 40384
rect 30929 40375 30987 40381
rect 30929 40372 30941 40375
rect 30800 40344 30941 40372
rect 30800 40332 30806 40344
rect 30929 40341 30941 40344
rect 30975 40341 30987 40375
rect 35342 40372 35348 40384
rect 35303 40344 35348 40372
rect 30929 40335 30987 40341
rect 35342 40332 35348 40344
rect 35400 40332 35406 40384
rect 36354 40372 36360 40384
rect 36315 40344 36360 40372
rect 36354 40332 36360 40344
rect 36412 40332 36418 40384
rect 36538 40332 36544 40384
rect 36596 40372 36602 40384
rect 37185 40375 37243 40381
rect 37185 40372 37197 40375
rect 36596 40344 37197 40372
rect 36596 40332 36602 40344
rect 37185 40341 37197 40344
rect 37231 40341 37243 40375
rect 37185 40335 37243 40341
rect 37277 40375 37335 40381
rect 37277 40341 37289 40375
rect 37323 40372 37335 40375
rect 37458 40372 37464 40384
rect 37323 40344 37464 40372
rect 37323 40341 37335 40344
rect 37277 40335 37335 40341
rect 37458 40332 37464 40344
rect 37516 40372 37522 40384
rect 41230 40372 41236 40384
rect 37516 40344 41236 40372
rect 37516 40332 37522 40344
rect 41230 40332 41236 40344
rect 41288 40332 41294 40384
rect 42518 40372 42524 40384
rect 42479 40344 42524 40372
rect 42518 40332 42524 40344
rect 42576 40332 42582 40384
rect 42978 40332 42984 40384
rect 43036 40372 43042 40384
rect 43349 40375 43407 40381
rect 43349 40372 43361 40375
rect 43036 40344 43361 40372
rect 43036 40332 43042 40344
rect 43349 40341 43361 40344
rect 43395 40341 43407 40375
rect 44174 40372 44180 40384
rect 44135 40344 44180 40372
rect 43349 40335 43407 40341
rect 44174 40332 44180 40344
rect 44232 40332 44238 40384
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 23842 40128 23848 40180
rect 23900 40168 23906 40180
rect 25869 40171 25927 40177
rect 23900 40140 24900 40168
rect 23900 40128 23906 40140
rect 23474 40060 23480 40112
rect 23532 40100 23538 40112
rect 23532 40072 23888 40100
rect 23532 40060 23538 40072
rect 23860 40041 23888 40072
rect 24394 40060 24400 40112
rect 24452 40100 24458 40112
rect 24734 40103 24792 40109
rect 24734 40100 24746 40103
rect 24452 40072 24746 40100
rect 24452 40060 24458 40072
rect 24734 40069 24746 40072
rect 24780 40069 24792 40103
rect 24872 40100 24900 40140
rect 25869 40137 25881 40171
rect 25915 40168 25927 40171
rect 27982 40168 27988 40180
rect 25915 40140 27988 40168
rect 25915 40137 25927 40140
rect 25869 40131 25927 40137
rect 27982 40128 27988 40140
rect 28040 40128 28046 40180
rect 35894 40128 35900 40180
rect 35952 40168 35958 40180
rect 37550 40168 37556 40180
rect 35952 40140 37556 40168
rect 35952 40128 35958 40140
rect 37550 40128 37556 40140
rect 37608 40128 37614 40180
rect 43901 40171 43959 40177
rect 43901 40137 43913 40171
rect 43947 40168 43959 40171
rect 44082 40168 44088 40180
rect 43947 40140 44088 40168
rect 43947 40137 43959 40140
rect 43901 40131 43959 40137
rect 44082 40128 44088 40140
rect 44140 40128 44146 40180
rect 44726 40128 44732 40180
rect 44784 40168 44790 40180
rect 46385 40171 46443 40177
rect 46385 40168 46397 40171
rect 44784 40140 46397 40168
rect 44784 40128 44790 40140
rect 46385 40137 46397 40140
rect 46431 40137 46443 40171
rect 46385 40131 46443 40137
rect 27246 40100 27252 40112
rect 24872 40072 27252 40100
rect 24734 40063 24792 40069
rect 27246 40060 27252 40072
rect 27304 40060 27310 40112
rect 29546 40100 29552 40112
rect 27356 40072 29552 40100
rect 23845 40035 23903 40041
rect 23845 40001 23857 40035
rect 23891 40001 23903 40035
rect 27157 40035 27215 40041
rect 27157 40032 27169 40035
rect 23845 39995 23903 40001
rect 25516 40004 27169 40032
rect 24489 39967 24547 39973
rect 24489 39933 24501 39967
rect 24535 39933 24547 39967
rect 24489 39927 24547 39933
rect 23658 39828 23664 39840
rect 23619 39800 23664 39828
rect 23658 39788 23664 39800
rect 23716 39788 23722 39840
rect 24504 39828 24532 39927
rect 24854 39828 24860 39840
rect 24504 39800 24860 39828
rect 24854 39788 24860 39800
rect 24912 39828 24918 39840
rect 25516 39828 25544 40004
rect 27157 40001 27169 40004
rect 27203 40032 27215 40035
rect 27356 40032 27384 40072
rect 29546 40060 29552 40072
rect 29604 40060 29610 40112
rect 44174 40100 44180 40112
rect 44100 40072 44180 40100
rect 27203 40004 27384 40032
rect 27424 40035 27482 40041
rect 27203 40001 27215 40004
rect 27157 39995 27215 40001
rect 27424 40001 27436 40035
rect 27470 40032 27482 40035
rect 29178 40032 29184 40044
rect 27470 40004 28212 40032
rect 29139 40004 29184 40032
rect 27470 40001 27482 40004
rect 27424 39995 27482 40001
rect 28184 39896 28212 40004
rect 29178 39992 29184 40004
rect 29236 39992 29242 40044
rect 30190 40032 30196 40044
rect 30103 40004 30196 40032
rect 30190 39992 30196 40004
rect 30248 40032 30254 40044
rect 31754 40032 31760 40044
rect 30248 40004 31760 40032
rect 30248 39992 30254 40004
rect 31754 39992 31760 40004
rect 31812 39992 31818 40044
rect 44100 40041 44128 40072
rect 44174 40060 44180 40072
rect 44232 40060 44238 40112
rect 44085 40035 44143 40041
rect 44085 40001 44097 40035
rect 44131 40001 44143 40035
rect 44085 39995 44143 40001
rect 45272 40035 45330 40041
rect 45272 40001 45284 40035
rect 45318 40032 45330 40035
rect 45830 40032 45836 40044
rect 45318 40004 45836 40032
rect 45318 40001 45330 40004
rect 45272 39995 45330 40001
rect 45830 39992 45836 40004
rect 45888 39992 45894 40044
rect 46845 40035 46903 40041
rect 46845 40001 46857 40035
rect 46891 40001 46903 40035
rect 46845 39995 46903 40001
rect 43990 39924 43996 39976
rect 44048 39964 44054 39976
rect 45005 39967 45063 39973
rect 45005 39964 45017 39967
rect 44048 39936 45017 39964
rect 44048 39924 44054 39936
rect 45005 39933 45017 39936
rect 45051 39933 45063 39967
rect 45005 39927 45063 39933
rect 28997 39899 29055 39905
rect 28997 39896 29009 39899
rect 28184 39868 29009 39896
rect 28997 39865 29009 39868
rect 29043 39865 29055 39899
rect 28997 39859 29055 39865
rect 31018 39856 31024 39908
rect 31076 39896 31082 39908
rect 46860 39896 46888 39995
rect 46934 39992 46940 40044
rect 46992 40032 46998 40044
rect 46992 40004 47037 40032
rect 46992 39992 46998 40004
rect 31076 39868 44128 39896
rect 31076 39856 31082 39868
rect 24912 39800 25544 39828
rect 24912 39788 24918 39800
rect 27890 39788 27896 39840
rect 27948 39828 27954 39840
rect 28537 39831 28595 39837
rect 28537 39828 28549 39831
rect 27948 39800 28549 39828
rect 27948 39788 27954 39800
rect 28537 39797 28549 39800
rect 28583 39797 28595 39831
rect 30006 39828 30012 39840
rect 29967 39800 30012 39828
rect 28537 39791 28595 39797
rect 30006 39788 30012 39800
rect 30064 39788 30070 39840
rect 44100 39828 44128 39868
rect 45940 39868 46888 39896
rect 45940 39828 45968 39868
rect 47762 39828 47768 39840
rect 44100 39800 45968 39828
rect 47723 39800 47768 39828
rect 47762 39788 47768 39800
rect 47820 39788 47826 39840
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 26602 39624 26608 39636
rect 26563 39596 26608 39624
rect 26602 39584 26608 39596
rect 26660 39584 26666 39636
rect 27062 39584 27068 39636
rect 27120 39624 27126 39636
rect 28629 39627 28687 39633
rect 28629 39624 28641 39627
rect 27120 39596 28641 39624
rect 27120 39584 27126 39596
rect 28629 39593 28641 39596
rect 28675 39593 28687 39627
rect 32582 39624 32588 39636
rect 32543 39596 32588 39624
rect 28629 39587 28687 39593
rect 32582 39584 32588 39596
rect 32640 39624 32646 39636
rect 38562 39624 38568 39636
rect 32640 39596 38568 39624
rect 32640 39584 32646 39596
rect 38562 39584 38568 39596
rect 38620 39624 38626 39636
rect 45094 39624 45100 39636
rect 38620 39596 45100 39624
rect 38620 39584 38626 39596
rect 45094 39584 45100 39596
rect 45152 39584 45158 39636
rect 27617 39559 27675 39565
rect 27617 39525 27629 39559
rect 27663 39556 27675 39559
rect 27982 39556 27988 39568
rect 27663 39528 27988 39556
rect 27663 39525 27675 39528
rect 27617 39519 27675 39525
rect 26237 39491 26295 39497
rect 26237 39457 26249 39491
rect 26283 39488 26295 39491
rect 27632 39488 27660 39519
rect 27982 39516 27988 39528
rect 28040 39516 28046 39568
rect 36630 39556 36636 39568
rect 32416 39528 36636 39556
rect 26283 39460 27660 39488
rect 26283 39457 26295 39460
rect 26237 39451 26295 39457
rect 24397 39423 24455 39429
rect 24397 39389 24409 39423
rect 24443 39420 24455 39423
rect 26421 39423 26479 39429
rect 24443 39392 24900 39420
rect 24443 39389 24455 39392
rect 24397 39383 24455 39389
rect 24872 39364 24900 39392
rect 26421 39389 26433 39423
rect 26467 39420 26479 39423
rect 27062 39420 27068 39432
rect 26467 39392 27068 39420
rect 26467 39389 26479 39392
rect 26421 39383 26479 39389
rect 27062 39380 27068 39392
rect 27120 39380 27126 39432
rect 27890 39420 27896 39432
rect 27851 39392 27896 39420
rect 27890 39380 27896 39392
rect 27948 39380 27954 39432
rect 28813 39423 28871 39429
rect 28813 39389 28825 39423
rect 28859 39420 28871 39423
rect 30190 39420 30196 39432
rect 28859 39392 30196 39420
rect 28859 39389 28871 39392
rect 28813 39383 28871 39389
rect 30190 39380 30196 39392
rect 30248 39380 30254 39432
rect 30742 39420 30748 39432
rect 30703 39392 30748 39420
rect 30742 39380 30748 39392
rect 30800 39380 30806 39432
rect 30834 39380 30840 39432
rect 30892 39420 30898 39432
rect 31021 39423 31079 39429
rect 30892 39392 30937 39420
rect 30892 39380 30898 39392
rect 31021 39389 31033 39423
rect 31067 39420 31079 39423
rect 31665 39423 31723 39429
rect 31665 39420 31677 39423
rect 31067 39392 31677 39420
rect 31067 39389 31079 39392
rect 31021 39383 31079 39389
rect 31665 39389 31677 39392
rect 31711 39389 31723 39423
rect 31665 39383 31723 39389
rect 31754 39380 31760 39432
rect 31812 39420 31818 39432
rect 32416 39429 32444 39528
rect 36630 39516 36636 39528
rect 36688 39516 36694 39568
rect 35894 39488 35900 39500
rect 35084 39460 35900 39488
rect 32401 39423 32459 39429
rect 32401 39420 32413 39423
rect 31812 39392 32413 39420
rect 31812 39380 31818 39392
rect 32401 39389 32413 39392
rect 32447 39389 32459 39423
rect 32401 39383 32459 39389
rect 34790 39380 34796 39432
rect 34848 39420 34854 39432
rect 35084 39429 35112 39460
rect 35894 39448 35900 39460
rect 35952 39448 35958 39500
rect 39114 39448 39120 39500
rect 39172 39488 39178 39500
rect 42794 39488 42800 39500
rect 39172 39460 42800 39488
rect 39172 39448 39178 39460
rect 42794 39448 42800 39460
rect 42852 39448 42858 39500
rect 46293 39491 46351 39497
rect 46293 39457 46305 39491
rect 46339 39488 46351 39491
rect 47762 39488 47768 39500
rect 46339 39460 47768 39488
rect 46339 39457 46351 39460
rect 46293 39451 46351 39457
rect 47762 39448 47768 39460
rect 47820 39448 47826 39500
rect 35342 39429 35348 39432
rect 34977 39423 35035 39429
rect 34977 39420 34989 39423
rect 34848 39392 34989 39420
rect 34848 39380 34854 39392
rect 34977 39389 34989 39392
rect 35023 39389 35035 39423
rect 34977 39383 35035 39389
rect 35069 39423 35127 39429
rect 35069 39389 35081 39423
rect 35115 39389 35127 39423
rect 35069 39383 35127 39389
rect 35299 39423 35348 39429
rect 35299 39389 35311 39423
rect 35345 39389 35348 39423
rect 35299 39383 35348 39389
rect 35342 39380 35348 39383
rect 35400 39380 35406 39432
rect 35434 39380 35440 39432
rect 35492 39420 35498 39432
rect 41877 39423 41935 39429
rect 35492 39392 35537 39420
rect 35492 39380 35498 39392
rect 41877 39389 41889 39423
rect 41923 39420 41935 39423
rect 42518 39420 42524 39432
rect 41923 39392 42524 39420
rect 41923 39389 41935 39392
rect 41877 39383 41935 39389
rect 42518 39380 42524 39392
rect 42576 39380 42582 39432
rect 42978 39420 42984 39432
rect 42939 39392 42984 39420
rect 42978 39380 42984 39392
rect 43036 39380 43042 39432
rect 23658 39312 23664 39364
rect 23716 39352 23722 39364
rect 24642 39355 24700 39361
rect 24642 39352 24654 39355
rect 23716 39324 24654 39352
rect 23716 39312 23722 39324
rect 24642 39321 24654 39324
rect 24688 39321 24700 39355
rect 24642 39315 24700 39321
rect 24854 39312 24860 39364
rect 24912 39312 24918 39364
rect 27706 39312 27712 39364
rect 27764 39352 27770 39364
rect 27985 39355 28043 39361
rect 27985 39352 27997 39355
rect 27764 39324 27997 39352
rect 27764 39312 27770 39324
rect 27985 39321 27997 39324
rect 28031 39321 28043 39355
rect 27985 39315 28043 39321
rect 35161 39355 35219 39361
rect 35161 39321 35173 39355
rect 35207 39352 35219 39355
rect 39298 39352 39304 39364
rect 35207 39324 39304 39352
rect 35207 39321 35219 39324
rect 35161 39315 35219 39321
rect 39298 39312 39304 39324
rect 39356 39312 39362 39364
rect 40402 39312 40408 39364
rect 40460 39352 40466 39364
rect 41693 39355 41751 39361
rect 40460 39324 41414 39352
rect 40460 39312 40466 39324
rect 25682 39244 25688 39296
rect 25740 39284 25746 39296
rect 25777 39287 25835 39293
rect 25777 39284 25789 39287
rect 25740 39256 25789 39284
rect 25740 39244 25746 39256
rect 25777 39253 25789 39256
rect 25823 39253 25835 39287
rect 27798 39284 27804 39296
rect 27759 39256 27804 39284
rect 25777 39247 25835 39253
rect 27798 39244 27804 39256
rect 27856 39244 27862 39296
rect 28169 39287 28227 39293
rect 28169 39253 28181 39287
rect 28215 39284 28227 39287
rect 28534 39284 28540 39296
rect 28215 39256 28540 39284
rect 28215 39253 28227 39256
rect 28169 39247 28227 39253
rect 28534 39244 28540 39256
rect 28592 39244 28598 39296
rect 31478 39284 31484 39296
rect 31439 39256 31484 39284
rect 31478 39244 31484 39256
rect 31536 39244 31542 39296
rect 34790 39284 34796 39296
rect 34751 39256 34796 39284
rect 34790 39244 34796 39256
rect 34848 39244 34854 39296
rect 41386 39284 41414 39324
rect 41693 39321 41705 39355
rect 41739 39352 41751 39355
rect 42334 39352 42340 39364
rect 41739 39324 42340 39352
rect 41739 39321 41751 39324
rect 41693 39315 41751 39321
rect 42334 39312 42340 39324
rect 42392 39312 42398 39364
rect 46477 39355 46535 39361
rect 46477 39321 46489 39355
rect 46523 39352 46535 39355
rect 47670 39352 47676 39364
rect 46523 39324 47676 39352
rect 46523 39321 46535 39324
rect 46477 39315 46535 39321
rect 47670 39312 47676 39324
rect 47728 39312 47734 39364
rect 48130 39352 48136 39364
rect 48091 39324 48136 39352
rect 48130 39312 48136 39324
rect 48188 39312 48194 39364
rect 42061 39287 42119 39293
rect 42061 39284 42073 39287
rect 41386 39256 42073 39284
rect 42061 39253 42073 39256
rect 42107 39253 42119 39287
rect 42061 39247 42119 39253
rect 42702 39244 42708 39296
rect 42760 39284 42766 39296
rect 42797 39287 42855 39293
rect 42797 39284 42809 39287
rect 42760 39256 42809 39284
rect 42760 39244 42766 39256
rect 42797 39253 42809 39256
rect 42843 39253 42855 39287
rect 42797 39247 42855 39253
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 24578 39040 24584 39092
rect 24636 39080 24642 39092
rect 31018 39080 31024 39092
rect 24636 39052 31024 39080
rect 24636 39040 24642 39052
rect 31018 39040 31024 39052
rect 31076 39040 31082 39092
rect 35434 39040 35440 39092
rect 35492 39080 35498 39092
rect 36357 39083 36415 39089
rect 36357 39080 36369 39083
rect 35492 39052 36369 39080
rect 35492 39040 35498 39052
rect 36357 39049 36369 39052
rect 36403 39049 36415 39083
rect 41046 39080 41052 39092
rect 36357 39043 36415 39049
rect 39224 39052 40540 39080
rect 41007 39052 41052 39080
rect 30834 38972 30840 39024
rect 30892 39012 30898 39024
rect 30892 38984 31754 39012
rect 30892 38972 30898 38984
rect 30006 38944 30012 38956
rect 29919 38916 30012 38944
rect 30006 38904 30012 38916
rect 30064 38944 30070 38956
rect 30852 38944 30880 38972
rect 30064 38916 30880 38944
rect 31726 38944 31754 38984
rect 31846 38972 31852 39024
rect 31904 39012 31910 39024
rect 33956 39015 34014 39021
rect 31904 38984 32444 39012
rect 31904 38972 31910 38984
rect 32309 38947 32367 38953
rect 32309 38944 32321 38947
rect 31726 38916 32321 38944
rect 30064 38904 30070 38916
rect 32309 38913 32321 38916
rect 32355 38913 32367 38947
rect 32416 38944 32444 38984
rect 33956 38981 33968 39015
rect 34002 39012 34014 39015
rect 35452 39012 35480 39040
rect 39224 39021 39252 39052
rect 39209 39015 39267 39021
rect 34002 38984 35480 39012
rect 35728 38984 37596 39012
rect 34002 38981 34014 38984
rect 33956 38975 34014 38981
rect 35728 38953 35756 38984
rect 37568 38953 37596 38984
rect 39209 38981 39221 39015
rect 39255 38981 39267 39015
rect 39209 38975 39267 38981
rect 39439 39015 39497 39021
rect 39439 38981 39451 39015
rect 39485 39012 39497 39015
rect 40402 39012 40408 39024
rect 39485 38984 40408 39012
rect 39485 38981 39497 38984
rect 39439 38975 39497 38981
rect 40402 38972 40408 38984
rect 40460 38972 40466 39024
rect 35713 38947 35771 38953
rect 35713 38944 35725 38947
rect 32416 38916 35725 38944
rect 32309 38907 32367 38913
rect 35713 38913 35725 38916
rect 35759 38913 35771 38947
rect 35713 38907 35771 38913
rect 35897 38947 35955 38953
rect 35897 38913 35909 38947
rect 35943 38944 35955 38947
rect 36541 38947 36599 38953
rect 36541 38944 36553 38947
rect 35943 38916 36553 38944
rect 35943 38913 35955 38916
rect 35897 38907 35955 38913
rect 36541 38913 36553 38916
rect 36587 38913 36599 38947
rect 36541 38907 36599 38913
rect 37553 38947 37611 38953
rect 37553 38913 37565 38947
rect 37599 38913 37611 38947
rect 37553 38907 37611 38913
rect 37737 38947 37795 38953
rect 37737 38913 37749 38947
rect 37783 38944 37795 38947
rect 38381 38947 38439 38953
rect 38381 38944 38393 38947
rect 37783 38916 38393 38944
rect 37783 38913 37795 38916
rect 37737 38907 37795 38913
rect 38381 38913 38393 38916
rect 38427 38913 38439 38947
rect 39114 38944 39120 38956
rect 39075 38916 39120 38944
rect 38381 38907 38439 38913
rect 29825 38879 29883 38885
rect 29825 38845 29837 38879
rect 29871 38876 29883 38879
rect 30190 38876 30196 38888
rect 29871 38848 30196 38876
rect 29871 38845 29883 38848
rect 29825 38839 29883 38845
rect 30190 38836 30196 38848
rect 30248 38836 30254 38888
rect 30745 38879 30803 38885
rect 30745 38845 30757 38879
rect 30791 38876 30803 38879
rect 30926 38876 30932 38888
rect 30791 38848 30932 38876
rect 30791 38845 30803 38848
rect 30745 38839 30803 38845
rect 30926 38836 30932 38848
rect 30984 38836 30990 38888
rect 31021 38879 31079 38885
rect 31021 38845 31033 38879
rect 31067 38876 31079 38879
rect 31754 38876 31760 38888
rect 31067 38848 31760 38876
rect 31067 38845 31079 38848
rect 31021 38839 31079 38845
rect 31754 38836 31760 38848
rect 31812 38836 31818 38888
rect 32125 38879 32183 38885
rect 32125 38845 32137 38879
rect 32171 38876 32183 38879
rect 32214 38876 32220 38888
rect 32171 38848 32220 38876
rect 32171 38845 32183 38848
rect 32125 38839 32183 38845
rect 32214 38836 32220 38848
rect 32272 38836 32278 38888
rect 33686 38876 33692 38888
rect 33647 38848 33692 38876
rect 33686 38836 33692 38848
rect 33744 38836 33750 38888
rect 35342 38836 35348 38888
rect 35400 38876 35406 38888
rect 35529 38879 35587 38885
rect 35529 38876 35541 38879
rect 35400 38848 35541 38876
rect 35400 38836 35406 38848
rect 35529 38845 35541 38848
rect 35575 38845 35587 38879
rect 35529 38839 35587 38845
rect 37090 38836 37096 38888
rect 37148 38876 37154 38888
rect 37369 38879 37427 38885
rect 37369 38876 37381 38879
rect 37148 38848 37381 38876
rect 37148 38836 37154 38848
rect 37369 38845 37381 38848
rect 37415 38845 37427 38879
rect 37568 38876 37596 38907
rect 39114 38904 39120 38916
rect 39172 38904 39178 38956
rect 39298 38904 39304 38956
rect 39356 38944 39362 38956
rect 40221 38947 40279 38953
rect 39356 38916 39712 38944
rect 39356 38904 39362 38916
rect 37826 38876 37832 38888
rect 37568 38848 37832 38876
rect 37369 38839 37427 38845
rect 37826 38836 37832 38848
rect 37884 38836 37890 38888
rect 39577 38879 39635 38885
rect 39577 38876 39589 38879
rect 38212 38848 39589 38876
rect 38212 38820 38240 38848
rect 39577 38845 39589 38848
rect 39623 38845 39635 38879
rect 39577 38839 39635 38845
rect 38194 38808 38200 38820
rect 38107 38780 38200 38808
rect 38194 38768 38200 38780
rect 38252 38768 38258 38820
rect 39684 38808 39712 38916
rect 40221 38913 40233 38947
rect 40267 38913 40279 38947
rect 40512 38944 40540 39052
rect 41046 39040 41052 39052
rect 41104 39040 41110 39092
rect 41141 39083 41199 39089
rect 41141 39049 41153 39083
rect 41187 39080 41199 39083
rect 41874 39080 41880 39092
rect 41187 39052 41880 39080
rect 41187 39049 41199 39052
rect 41141 39043 41199 39049
rect 41874 39040 41880 39052
rect 41932 39040 41938 39092
rect 47670 39080 47676 39092
rect 47631 39052 47676 39080
rect 47670 39040 47676 39052
rect 47728 39040 47734 39092
rect 40957 39015 41015 39021
rect 40957 38981 40969 39015
rect 41003 39012 41015 39015
rect 41414 39012 41420 39024
rect 41003 38984 41420 39012
rect 41003 38981 41015 38984
rect 40957 38975 41015 38981
rect 41414 38972 41420 38984
rect 41472 38972 41478 39024
rect 42444 38984 44036 39012
rect 42444 38953 42472 38984
rect 44008 38956 44036 38984
rect 42702 38953 42708 38956
rect 42429 38947 42487 38953
rect 40512 38916 41092 38944
rect 40221 38907 40279 38913
rect 40236 38876 40264 38907
rect 41064 38876 41092 38916
rect 42429 38913 42441 38947
rect 42475 38913 42487 38947
rect 42696 38944 42708 38953
rect 42663 38916 42708 38944
rect 42429 38907 42487 38913
rect 42696 38907 42708 38916
rect 42702 38904 42708 38907
rect 42760 38904 42766 38956
rect 43990 38904 43996 38956
rect 44048 38944 44054 38956
rect 45189 38947 45247 38953
rect 45189 38944 45201 38947
rect 44048 38916 45201 38944
rect 44048 38904 44054 38916
rect 45189 38913 45201 38916
rect 45235 38913 45247 38947
rect 45189 38907 45247 38913
rect 45456 38947 45514 38953
rect 45456 38913 45468 38947
rect 45502 38944 45514 38947
rect 46750 38944 46756 38956
rect 45502 38916 46756 38944
rect 45502 38913 45514 38916
rect 45456 38907 45514 38913
rect 41325 38879 41383 38885
rect 41325 38876 41337 38879
rect 40236 38848 41000 38876
rect 41064 38848 41337 38876
rect 40586 38808 40592 38820
rect 39684 38780 40592 38808
rect 40586 38768 40592 38780
rect 40644 38768 40650 38820
rect 40770 38808 40776 38820
rect 40731 38780 40776 38808
rect 40770 38768 40776 38780
rect 40828 38768 40834 38820
rect 40972 38808 41000 38848
rect 41325 38845 41337 38848
rect 41371 38845 41383 38879
rect 41325 38839 41383 38845
rect 41782 38808 41788 38820
rect 40972 38780 41788 38808
rect 41782 38768 41788 38780
rect 41840 38768 41846 38820
rect 29822 38700 29828 38752
rect 29880 38740 29886 38752
rect 30193 38743 30251 38749
rect 30193 38740 30205 38743
rect 29880 38712 30205 38740
rect 29880 38700 29886 38712
rect 30193 38709 30205 38712
rect 30239 38709 30251 38743
rect 30193 38703 30251 38709
rect 32493 38743 32551 38749
rect 32493 38709 32505 38743
rect 32539 38740 32551 38743
rect 32858 38740 32864 38752
rect 32539 38712 32864 38740
rect 32539 38709 32551 38712
rect 32493 38703 32551 38709
rect 32858 38700 32864 38712
rect 32916 38700 32922 38752
rect 35069 38743 35127 38749
rect 35069 38709 35081 38743
rect 35115 38740 35127 38743
rect 35618 38740 35624 38752
rect 35115 38712 35624 38740
rect 35115 38709 35127 38712
rect 35069 38703 35127 38709
rect 35618 38700 35624 38712
rect 35676 38700 35682 38752
rect 38930 38740 38936 38752
rect 38891 38712 38936 38740
rect 38930 38700 38936 38712
rect 38988 38700 38994 38752
rect 40037 38743 40095 38749
rect 40037 38709 40049 38743
rect 40083 38740 40095 38743
rect 40126 38740 40132 38752
rect 40083 38712 40132 38740
rect 40083 38709 40095 38712
rect 40037 38703 40095 38709
rect 40126 38700 40132 38712
rect 40184 38700 40190 38752
rect 41414 38700 41420 38752
rect 41472 38740 41478 38752
rect 42150 38740 42156 38752
rect 41472 38712 42156 38740
rect 41472 38700 41478 38712
rect 42150 38700 42156 38712
rect 42208 38740 42214 38752
rect 43809 38743 43867 38749
rect 43809 38740 43821 38743
rect 42208 38712 43821 38740
rect 42208 38700 42214 38712
rect 43809 38709 43821 38712
rect 43855 38709 43867 38743
rect 45204 38740 45232 38907
rect 46750 38904 46756 38916
rect 46808 38904 46814 38956
rect 47578 38944 47584 38956
rect 47539 38916 47584 38944
rect 47578 38904 47584 38916
rect 47636 38904 47642 38956
rect 45554 38740 45560 38752
rect 45204 38712 45560 38740
rect 43809 38703 43867 38709
rect 45554 38700 45560 38712
rect 45612 38700 45618 38752
rect 46566 38740 46572 38752
rect 46527 38712 46572 38740
rect 46566 38700 46572 38712
rect 46624 38700 46630 38752
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 26050 38496 26056 38548
rect 26108 38536 26114 38548
rect 40954 38536 40960 38548
rect 26108 38508 40960 38536
rect 26108 38496 26114 38508
rect 40954 38496 40960 38508
rect 41012 38496 41018 38548
rect 41046 38496 41052 38548
rect 41104 38536 41110 38548
rect 41598 38536 41604 38548
rect 41104 38508 41604 38536
rect 41104 38496 41110 38508
rect 41598 38496 41604 38508
rect 41656 38496 41662 38548
rect 42058 38496 42064 38548
rect 42116 38536 42122 38548
rect 42334 38536 42340 38548
rect 42116 38508 42161 38536
rect 42295 38508 42340 38536
rect 42116 38496 42122 38508
rect 42334 38496 42340 38508
rect 42392 38496 42398 38548
rect 46750 38536 46756 38548
rect 46711 38508 46756 38536
rect 46750 38496 46756 38508
rect 46808 38496 46814 38548
rect 32214 38468 32220 38480
rect 32175 38440 32220 38468
rect 32214 38428 32220 38440
rect 32272 38428 32278 38480
rect 29546 38360 29552 38412
rect 29604 38400 29610 38412
rect 30377 38403 30435 38409
rect 30377 38400 30389 38403
rect 29604 38372 30389 38400
rect 29604 38360 29610 38372
rect 30377 38369 30389 38372
rect 30423 38369 30435 38403
rect 33686 38400 33692 38412
rect 30377 38363 30435 38369
rect 32140 38372 33692 38400
rect 32140 38344 32168 38372
rect 33686 38360 33692 38372
rect 33744 38400 33750 38412
rect 34701 38403 34759 38409
rect 34701 38400 34713 38403
rect 33744 38372 34713 38400
rect 33744 38360 33750 38372
rect 34701 38369 34713 38372
rect 34747 38369 34759 38403
rect 34701 38363 34759 38369
rect 42058 38360 42064 38412
rect 42116 38400 42122 38412
rect 45922 38400 45928 38412
rect 42116 38372 42161 38400
rect 45835 38372 45928 38400
rect 42116 38360 42122 38372
rect 45922 38360 45928 38372
rect 45980 38400 45986 38412
rect 46566 38400 46572 38412
rect 45980 38372 46572 38400
rect 45980 38360 45986 38372
rect 46566 38360 46572 38372
rect 46624 38360 46630 38412
rect 25774 38332 25780 38344
rect 25735 38304 25780 38332
rect 25774 38292 25780 38304
rect 25832 38292 25838 38344
rect 28166 38292 28172 38344
rect 28224 38332 28230 38344
rect 28721 38335 28779 38341
rect 28721 38332 28733 38335
rect 28224 38304 28733 38332
rect 28224 38292 28230 38304
rect 28721 38301 28733 38304
rect 28767 38301 28779 38335
rect 28721 38295 28779 38301
rect 30009 38335 30067 38341
rect 30009 38301 30021 38335
rect 30055 38332 30067 38335
rect 30742 38332 30748 38344
rect 30055 38304 30748 38332
rect 30055 38301 30067 38304
rect 30009 38295 30067 38301
rect 30742 38292 30748 38304
rect 30800 38292 30806 38344
rect 30837 38335 30895 38341
rect 30837 38301 30849 38335
rect 30883 38332 30895 38335
rect 32122 38332 32128 38344
rect 30883 38304 32128 38332
rect 30883 38301 30895 38304
rect 30837 38295 30895 38301
rect 32122 38292 32128 38304
rect 32180 38292 32186 38344
rect 32858 38332 32864 38344
rect 32819 38304 32864 38332
rect 32858 38292 32864 38304
rect 32916 38292 32922 38344
rect 34790 38292 34796 38344
rect 34848 38332 34854 38344
rect 34957 38335 35015 38341
rect 34957 38332 34969 38335
rect 34848 38304 34969 38332
rect 34848 38292 34854 38304
rect 34957 38301 34969 38304
rect 35003 38301 35015 38335
rect 37182 38332 37188 38344
rect 37143 38304 37188 38332
rect 34957 38295 35015 38301
rect 37182 38292 37188 38304
rect 37240 38292 37246 38344
rect 37452 38335 37510 38341
rect 37452 38301 37464 38335
rect 37498 38332 37510 38335
rect 38194 38332 38200 38344
rect 37498 38304 38200 38332
rect 37498 38301 37510 38304
rect 37452 38295 37510 38301
rect 38194 38292 38200 38304
rect 38252 38292 38258 38344
rect 40037 38335 40095 38341
rect 40037 38301 40049 38335
rect 40083 38301 40095 38335
rect 40037 38295 40095 38301
rect 28537 38267 28595 38273
rect 28537 38233 28549 38267
rect 28583 38264 28595 38267
rect 29730 38264 29736 38276
rect 28583 38236 29736 38264
rect 28583 38233 28595 38236
rect 28537 38227 28595 38233
rect 29730 38224 29736 38236
rect 29788 38224 29794 38276
rect 29825 38267 29883 38273
rect 29825 38233 29837 38267
rect 29871 38264 29883 38267
rect 31104 38267 31162 38273
rect 29871 38236 31064 38264
rect 29871 38233 29883 38236
rect 29825 38227 29883 38233
rect 25590 38196 25596 38208
rect 25551 38168 25596 38196
rect 25590 38156 25596 38168
rect 25648 38156 25654 38208
rect 28902 38196 28908 38208
rect 28863 38168 28908 38196
rect 28902 38156 28908 38168
rect 28960 38156 28966 38208
rect 30098 38196 30104 38208
rect 30059 38168 30104 38196
rect 30098 38156 30104 38168
rect 30156 38156 30162 38208
rect 30190 38156 30196 38208
rect 30248 38196 30254 38208
rect 31036 38196 31064 38236
rect 31104 38233 31116 38267
rect 31150 38264 31162 38267
rect 31478 38264 31484 38276
rect 31150 38236 31484 38264
rect 31150 38233 31162 38236
rect 31104 38227 31162 38233
rect 31478 38224 31484 38236
rect 31536 38224 31542 38276
rect 31294 38196 31300 38208
rect 30248 38168 30293 38196
rect 31036 38168 31300 38196
rect 30248 38156 30254 38168
rect 31294 38156 31300 38168
rect 31352 38196 31358 38208
rect 32214 38196 32220 38208
rect 31352 38168 32220 38196
rect 31352 38156 31358 38168
rect 32214 38156 32220 38168
rect 32272 38156 32278 38208
rect 32674 38196 32680 38208
rect 32635 38168 32680 38196
rect 32674 38156 32680 38168
rect 32732 38156 32738 38208
rect 35342 38156 35348 38208
rect 35400 38196 35406 38208
rect 36081 38199 36139 38205
rect 36081 38196 36093 38199
rect 35400 38168 36093 38196
rect 35400 38156 35406 38168
rect 36081 38165 36093 38168
rect 36127 38165 36139 38199
rect 36081 38159 36139 38165
rect 36446 38156 36452 38208
rect 36504 38196 36510 38208
rect 38565 38199 38623 38205
rect 38565 38196 38577 38199
rect 36504 38168 38577 38196
rect 36504 38156 36510 38168
rect 38565 38165 38577 38168
rect 38611 38165 38623 38199
rect 40052 38196 40080 38295
rect 40770 38292 40776 38344
rect 40828 38332 40834 38344
rect 42153 38335 42211 38341
rect 42153 38332 42165 38335
rect 40828 38304 42165 38332
rect 40828 38292 40834 38304
rect 42153 38301 42165 38304
rect 42199 38301 42211 38335
rect 42153 38295 42211 38301
rect 42794 38292 42800 38344
rect 42852 38332 42858 38344
rect 43073 38335 43131 38341
rect 43073 38332 43085 38335
rect 42852 38304 43085 38332
rect 42852 38292 42858 38304
rect 43073 38301 43085 38304
rect 43119 38332 43131 38335
rect 43898 38332 43904 38344
rect 43119 38304 43904 38332
rect 43119 38301 43131 38304
rect 43073 38295 43131 38301
rect 43898 38292 43904 38304
rect 43956 38292 43962 38344
rect 45094 38332 45100 38344
rect 45055 38304 45100 38332
rect 45094 38292 45100 38304
rect 45152 38292 45158 38344
rect 45189 38335 45247 38341
rect 45189 38301 45201 38335
rect 45235 38332 45247 38335
rect 46109 38335 46167 38341
rect 46109 38332 46121 38335
rect 45235 38304 46121 38332
rect 45235 38301 45247 38304
rect 45189 38295 45247 38301
rect 46109 38301 46121 38304
rect 46155 38301 46167 38335
rect 46109 38295 46167 38301
rect 46937 38335 46995 38341
rect 46937 38301 46949 38335
rect 46983 38301 46995 38335
rect 47394 38332 47400 38344
rect 47355 38304 47400 38332
rect 46937 38295 46995 38301
rect 40304 38267 40362 38273
rect 40304 38233 40316 38267
rect 40350 38264 40362 38267
rect 41506 38264 41512 38276
rect 40350 38236 41512 38264
rect 40350 38233 40362 38236
rect 40304 38227 40362 38233
rect 41506 38224 41512 38236
rect 41564 38224 41570 38276
rect 41874 38264 41880 38276
rect 41835 38236 41880 38264
rect 41874 38224 41880 38236
rect 41932 38224 41938 38276
rect 43340 38267 43398 38273
rect 43340 38233 43352 38267
rect 43386 38264 43398 38267
rect 43806 38264 43812 38276
rect 43386 38236 43812 38264
rect 43386 38233 43398 38236
rect 43340 38227 43398 38233
rect 43806 38224 43812 38236
rect 43864 38224 43870 38276
rect 44082 38224 44088 38276
rect 44140 38264 44146 38276
rect 45204 38264 45232 38295
rect 44140 38236 45232 38264
rect 45373 38267 45431 38273
rect 44140 38224 44146 38236
rect 45373 38233 45385 38267
rect 45419 38264 45431 38267
rect 46952 38264 46980 38295
rect 47394 38292 47400 38304
rect 47452 38292 47458 38344
rect 45419 38236 46980 38264
rect 45419 38233 45431 38236
rect 45373 38227 45431 38233
rect 40218 38196 40224 38208
rect 40052 38168 40224 38196
rect 38565 38159 38623 38165
rect 40218 38156 40224 38168
rect 40276 38196 40282 38208
rect 40494 38196 40500 38208
rect 40276 38168 40500 38196
rect 40276 38156 40282 38168
rect 40494 38156 40500 38168
rect 40552 38156 40558 38208
rect 41417 38199 41475 38205
rect 41417 38165 41429 38199
rect 41463 38196 41475 38199
rect 41598 38196 41604 38208
rect 41463 38168 41604 38196
rect 41463 38165 41475 38168
rect 41417 38159 41475 38165
rect 41598 38156 41604 38168
rect 41656 38196 41662 38208
rect 42058 38196 42064 38208
rect 41656 38168 42064 38196
rect 41656 38156 41662 38168
rect 42058 38156 42064 38168
rect 42116 38156 42122 38208
rect 44453 38199 44511 38205
rect 44453 38165 44465 38199
rect 44499 38196 44511 38199
rect 45094 38196 45100 38208
rect 44499 38168 45100 38196
rect 44499 38165 44511 38168
rect 44453 38159 44511 38165
rect 45094 38156 45100 38168
rect 45152 38156 45158 38208
rect 46290 38196 46296 38208
rect 46251 38168 46296 38196
rect 46290 38156 46296 38168
rect 46348 38156 46354 38208
rect 47486 38196 47492 38208
rect 47447 38168 47492 38196
rect 47486 38156 47492 38168
rect 47544 38156 47550 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 30098 37952 30104 38004
rect 30156 37992 30162 38004
rect 30561 37995 30619 38001
rect 30561 37992 30573 37995
rect 30156 37964 30573 37992
rect 30156 37952 30162 37964
rect 30561 37961 30573 37964
rect 30607 37992 30619 37995
rect 35618 37992 35624 38004
rect 30607 37964 31248 37992
rect 35579 37964 35624 37992
rect 30607 37961 30619 37964
rect 30561 37955 30619 37961
rect 27614 37924 27620 37936
rect 25056 37896 27620 37924
rect 24854 37748 24860 37800
rect 24912 37788 24918 37800
rect 25056 37797 25084 37896
rect 27614 37884 27620 37896
rect 27672 37924 27678 37936
rect 27672 37896 29224 37924
rect 27672 37884 27678 37896
rect 25308 37859 25366 37865
rect 25308 37825 25320 37859
rect 25354 37856 25366 37859
rect 25590 37856 25596 37868
rect 25354 37828 25596 37856
rect 25354 37825 25366 37828
rect 25308 37819 25366 37825
rect 25590 37816 25596 37828
rect 25648 37816 25654 37868
rect 29196 37865 29224 37896
rect 30190 37884 30196 37936
rect 30248 37924 30254 37936
rect 30248 37896 31064 37924
rect 30248 37884 30254 37896
rect 29454 37865 29460 37868
rect 29181 37859 29239 37865
rect 29181 37825 29193 37859
rect 29227 37825 29239 37859
rect 29181 37819 29239 37825
rect 29448 37819 29460 37865
rect 29512 37856 29518 37868
rect 29512 37828 29548 37856
rect 29454 37816 29460 37819
rect 29512 37816 29518 37828
rect 29730 37816 29736 37868
rect 29788 37856 29794 37868
rect 31036 37865 31064 37896
rect 31220 37865 31248 37964
rect 35618 37952 35624 37964
rect 35676 37952 35682 38004
rect 37090 37992 37096 38004
rect 35866 37964 37096 37992
rect 32392 37927 32450 37933
rect 32392 37893 32404 37927
rect 32438 37924 32450 37927
rect 32674 37924 32680 37936
rect 32438 37896 32680 37924
rect 32438 37893 32450 37896
rect 32392 37887 32450 37893
rect 32674 37884 32680 37896
rect 32732 37884 32738 37936
rect 35866 37933 35894 37964
rect 37090 37952 37096 37964
rect 37148 37992 37154 38004
rect 38657 37995 38715 38001
rect 38657 37992 38669 37995
rect 37148 37964 38669 37992
rect 37148 37952 37154 37964
rect 38657 37961 38669 37964
rect 38703 37961 38715 37995
rect 38657 37955 38715 37961
rect 40770 37952 40776 38004
rect 40828 37992 40834 38004
rect 40957 37995 41015 38001
rect 40957 37992 40969 37995
rect 40828 37964 40969 37992
rect 40828 37952 40834 37964
rect 40957 37961 40969 37964
rect 41003 37961 41015 37995
rect 41782 37992 41788 38004
rect 41743 37964 41788 37992
rect 40957 37955 41015 37961
rect 41782 37952 41788 37964
rect 41840 37952 41846 38004
rect 43806 37952 43812 38004
rect 43864 37992 43870 38004
rect 43901 37995 43959 38001
rect 43901 37992 43913 37995
rect 43864 37964 43913 37992
rect 43864 37952 43870 37964
rect 43901 37961 43913 37964
rect 43947 37961 43959 37995
rect 43901 37955 43959 37961
rect 47581 37995 47639 38001
rect 47581 37961 47593 37995
rect 47627 37961 47639 37995
rect 47581 37955 47639 37961
rect 35830 37927 35894 37933
rect 35830 37893 35842 37927
rect 35876 37896 35894 37927
rect 45916 37927 45974 37933
rect 35876 37893 35888 37896
rect 35830 37887 35888 37893
rect 45916 37893 45928 37927
rect 45962 37924 45974 37927
rect 47596 37924 47624 37955
rect 45962 37896 47624 37924
rect 45962 37893 45974 37896
rect 45916 37887 45974 37893
rect 31021 37859 31079 37865
rect 29788 37828 30236 37856
rect 29788 37816 29794 37828
rect 25041 37791 25099 37797
rect 25041 37788 25053 37791
rect 24912 37760 25053 37788
rect 24912 37748 24918 37760
rect 25041 37757 25053 37760
rect 25087 37757 25099 37791
rect 25041 37751 25099 37757
rect 30208 37720 30236 37828
rect 31021 37825 31033 37859
rect 31067 37825 31079 37859
rect 31021 37819 31079 37825
rect 31205 37859 31263 37865
rect 31205 37825 31217 37859
rect 31251 37825 31263 37859
rect 31205 37819 31263 37825
rect 31036 37788 31064 37819
rect 31294 37816 31300 37868
rect 31352 37856 31358 37868
rect 35710 37856 35716 37868
rect 31352 37828 31397 37856
rect 35623 37828 35716 37856
rect 31352 37816 31358 37828
rect 35710 37816 35716 37828
rect 35768 37856 35774 37868
rect 36446 37856 36452 37868
rect 35768 37828 36452 37856
rect 35768 37816 35774 37828
rect 36446 37816 36452 37828
rect 36504 37816 36510 37868
rect 36633 37859 36691 37865
rect 36633 37825 36645 37859
rect 36679 37825 36691 37859
rect 36633 37819 36691 37825
rect 32122 37788 32128 37800
rect 31036 37760 31616 37788
rect 32083 37760 32128 37788
rect 31481 37723 31539 37729
rect 31481 37720 31493 37723
rect 30208 37692 31493 37720
rect 31481 37689 31493 37692
rect 31527 37689 31539 37723
rect 31481 37683 31539 37689
rect 26421 37655 26479 37661
rect 26421 37621 26433 37655
rect 26467 37652 26479 37655
rect 26786 37652 26792 37664
rect 26467 37624 26792 37652
rect 26467 37621 26479 37624
rect 26421 37615 26479 37621
rect 26786 37612 26792 37624
rect 26844 37612 26850 37664
rect 30742 37612 30748 37664
rect 30800 37652 30806 37664
rect 31021 37655 31079 37661
rect 31021 37652 31033 37655
rect 30800 37624 31033 37652
rect 30800 37612 30806 37624
rect 31021 37621 31033 37624
rect 31067 37621 31079 37655
rect 31588 37652 31616 37760
rect 32122 37748 32128 37760
rect 32180 37748 32186 37800
rect 35342 37788 35348 37800
rect 35303 37760 35348 37788
rect 35342 37748 35348 37760
rect 35400 37748 35406 37800
rect 35618 37748 35624 37800
rect 35676 37788 35682 37800
rect 36648 37788 36676 37819
rect 37182 37816 37188 37868
rect 37240 37856 37246 37868
rect 37277 37859 37335 37865
rect 37277 37856 37289 37859
rect 37240 37828 37289 37856
rect 37240 37816 37246 37828
rect 37277 37825 37289 37828
rect 37323 37825 37335 37859
rect 37277 37819 37335 37825
rect 37544 37859 37602 37865
rect 37544 37825 37556 37859
rect 37590 37856 37602 37859
rect 38930 37856 38936 37868
rect 37590 37828 38936 37856
rect 37590 37825 37602 37828
rect 37544 37819 37602 37825
rect 35676 37760 36676 37788
rect 35676 37748 35682 37760
rect 33505 37655 33563 37661
rect 33505 37652 33517 37655
rect 31588 37624 33517 37652
rect 31021 37615 31079 37621
rect 33505 37621 33517 37624
rect 33551 37621 33563 37655
rect 35986 37652 35992 37664
rect 35947 37624 35992 37652
rect 33505 37615 33563 37621
rect 35986 37612 35992 37624
rect 36044 37612 36050 37664
rect 36262 37612 36268 37664
rect 36320 37652 36326 37664
rect 36449 37655 36507 37661
rect 36449 37652 36461 37655
rect 36320 37624 36461 37652
rect 36320 37612 36326 37624
rect 36449 37621 36461 37624
rect 36495 37621 36507 37655
rect 37292 37652 37320 37819
rect 38930 37816 38936 37828
rect 38988 37816 38994 37868
rect 39844 37859 39902 37865
rect 39844 37825 39856 37859
rect 39890 37856 39902 37859
rect 40126 37856 40132 37868
rect 39890 37828 40132 37856
rect 39890 37825 39902 37828
rect 39844 37819 39902 37825
rect 40126 37816 40132 37828
rect 40184 37816 40190 37868
rect 41414 37856 41420 37868
rect 41375 37828 41420 37856
rect 41414 37816 41420 37828
rect 41472 37816 41478 37868
rect 41601 37859 41659 37865
rect 41601 37825 41613 37859
rect 41647 37825 41659 37859
rect 41601 37819 41659 37825
rect 44085 37859 44143 37865
rect 44085 37825 44097 37859
rect 44131 37856 44143 37859
rect 44266 37856 44272 37868
rect 44131 37828 44272 37856
rect 44131 37825 44143 37828
rect 44085 37819 44143 37825
rect 39577 37791 39635 37797
rect 39577 37757 39589 37791
rect 39623 37757 39635 37791
rect 39577 37751 39635 37757
rect 39592 37652 39620 37751
rect 40954 37748 40960 37800
rect 41012 37788 41018 37800
rect 41616 37788 41644 37819
rect 44266 37816 44272 37828
rect 44324 37816 44330 37868
rect 45554 37816 45560 37868
rect 45612 37856 45618 37868
rect 45649 37859 45707 37865
rect 45649 37856 45661 37859
rect 45612 37828 45661 37856
rect 45612 37816 45618 37828
rect 45649 37825 45661 37828
rect 45695 37825 45707 37859
rect 45649 37819 45707 37825
rect 46290 37816 46296 37868
rect 46348 37856 46354 37868
rect 47765 37859 47823 37865
rect 47765 37856 47777 37859
rect 46348 37828 47777 37856
rect 46348 37816 46354 37828
rect 47765 37825 47777 37828
rect 47811 37825 47823 37859
rect 47765 37819 47823 37825
rect 41012 37760 41644 37788
rect 41012 37748 41018 37760
rect 40494 37652 40500 37664
rect 37292 37624 40500 37652
rect 36449 37615 36507 37621
rect 40494 37612 40500 37624
rect 40552 37612 40558 37664
rect 46934 37612 46940 37664
rect 46992 37652 46998 37664
rect 47029 37655 47087 37661
rect 47029 37652 47041 37655
rect 46992 37624 47041 37652
rect 46992 37612 46998 37624
rect 47029 37621 47041 37624
rect 47075 37621 47087 37655
rect 47029 37615 47087 37621
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 25774 37408 25780 37460
rect 25832 37448 25838 37460
rect 26145 37451 26203 37457
rect 26145 37448 26157 37451
rect 25832 37420 26157 37448
rect 25832 37408 25838 37420
rect 26145 37417 26157 37420
rect 26191 37417 26203 37451
rect 26145 37411 26203 37417
rect 29454 37408 29460 37460
rect 29512 37448 29518 37460
rect 29641 37451 29699 37457
rect 29641 37448 29653 37451
rect 29512 37420 29653 37448
rect 29512 37408 29518 37420
rect 29641 37417 29653 37420
rect 29687 37417 29699 37451
rect 41506 37448 41512 37460
rect 41467 37420 41512 37448
rect 29641 37411 29699 37417
rect 41506 37408 41512 37420
rect 41564 37408 41570 37460
rect 29546 37380 29552 37392
rect 28828 37352 29552 37380
rect 26786 37312 26792 37324
rect 26747 37284 26792 37312
rect 26786 37272 26792 37284
rect 26844 37312 26850 37324
rect 27062 37312 27068 37324
rect 26844 37284 27068 37312
rect 26844 37272 26850 37284
rect 27062 37272 27068 37284
rect 27120 37272 27126 37324
rect 28828 37312 28856 37352
rect 29546 37340 29552 37352
rect 29604 37340 29610 37392
rect 35618 37380 35624 37392
rect 34716 37352 35624 37380
rect 28994 37312 29000 37324
rect 28736 37284 28856 37312
rect 28955 37284 29000 37312
rect 24946 37244 24952 37256
rect 24907 37216 24952 37244
rect 24946 37204 24952 37216
rect 25004 37204 25010 37256
rect 25774 37244 25780 37256
rect 25735 37216 25780 37244
rect 25774 37204 25780 37216
rect 25832 37204 25838 37256
rect 25961 37247 26019 37253
rect 25961 37213 25973 37247
rect 26007 37244 26019 37247
rect 26970 37244 26976 37256
rect 26007 37216 26976 37244
rect 26007 37213 26019 37216
rect 25961 37207 26019 37213
rect 26970 37204 26976 37216
rect 27028 37204 27034 37256
rect 27157 37247 27215 37253
rect 27157 37213 27169 37247
rect 27203 37244 27215 37247
rect 27801 37247 27859 37253
rect 27801 37244 27813 37247
rect 27203 37216 27813 37244
rect 27203 37213 27215 37216
rect 27157 37207 27215 37213
rect 27801 37213 27813 37216
rect 27847 37213 27859 37247
rect 28534 37244 28540 37256
rect 28495 37216 28540 37244
rect 27801 37207 27859 37213
rect 28534 37204 28540 37216
rect 28592 37204 28598 37256
rect 28629 37247 28687 37253
rect 28629 37213 28641 37247
rect 28675 37244 28687 37247
rect 28736 37244 28764 37284
rect 28994 37272 29000 37284
rect 29052 37272 29058 37324
rect 34716 37321 34744 37352
rect 35618 37340 35624 37352
rect 35676 37340 35682 37392
rect 35805 37383 35863 37389
rect 35805 37349 35817 37383
rect 35851 37380 35863 37383
rect 36446 37380 36452 37392
rect 35851 37352 36452 37380
rect 35851 37349 35863 37352
rect 35805 37343 35863 37349
rect 36446 37340 36452 37352
rect 36504 37340 36510 37392
rect 36725 37383 36783 37389
rect 36725 37349 36737 37383
rect 36771 37349 36783 37383
rect 41874 37380 41880 37392
rect 36725 37343 36783 37349
rect 39868 37352 41880 37380
rect 34701 37315 34759 37321
rect 34701 37281 34713 37315
rect 34747 37281 34759 37315
rect 34701 37275 34759 37281
rect 35342 37272 35348 37324
rect 35400 37312 35406 37324
rect 35529 37315 35587 37321
rect 35529 37312 35541 37315
rect 35400 37284 35541 37312
rect 35400 37272 35406 37284
rect 35529 37281 35541 37284
rect 35575 37312 35587 37315
rect 36740 37312 36768 37343
rect 39868 37321 39896 37352
rect 41874 37340 41880 37352
rect 41932 37380 41938 37392
rect 42242 37380 42248 37392
rect 41932 37352 42248 37380
rect 41932 37340 41938 37352
rect 42242 37340 42248 37352
rect 42300 37340 42306 37392
rect 44082 37340 44088 37392
rect 44140 37340 44146 37392
rect 35575 37284 36768 37312
rect 39853 37315 39911 37321
rect 35575 37281 35587 37284
rect 35529 37275 35587 37281
rect 39853 37281 39865 37315
rect 39899 37281 39911 37315
rect 39853 37275 39911 37281
rect 40681 37315 40739 37321
rect 40681 37281 40693 37315
rect 40727 37312 40739 37315
rect 40770 37312 40776 37324
rect 40727 37284 40776 37312
rect 40727 37281 40739 37284
rect 40681 37275 40739 37281
rect 40770 37272 40776 37284
rect 40828 37272 40834 37324
rect 28902 37253 28908 37256
rect 28675 37216 28764 37244
rect 28859 37247 28908 37253
rect 28675 37213 28687 37216
rect 28629 37207 28687 37213
rect 28859 37213 28871 37247
rect 28905 37213 28908 37247
rect 28859 37207 28908 37213
rect 28902 37204 28908 37207
rect 28960 37204 28966 37256
rect 29822 37244 29828 37256
rect 29783 37216 29828 37244
rect 29822 37204 29828 37216
rect 29880 37204 29886 37256
rect 34885 37247 34943 37253
rect 34885 37213 34897 37247
rect 34931 37244 34943 37247
rect 35710 37244 35716 37256
rect 34931 37216 35716 37244
rect 34931 37213 34943 37216
rect 34885 37207 34943 37213
rect 35710 37204 35716 37216
rect 35768 37204 35774 37256
rect 36446 37244 36452 37256
rect 36359 37216 36452 37244
rect 36446 37204 36452 37216
rect 36504 37244 36510 37256
rect 37090 37244 37096 37256
rect 36504 37216 37096 37244
rect 36504 37204 36510 37216
rect 37090 37204 37096 37216
rect 37148 37204 37154 37256
rect 40037 37247 40095 37253
rect 40037 37213 40049 37247
rect 40083 37244 40095 37247
rect 40865 37247 40923 37253
rect 40865 37244 40877 37247
rect 40083 37216 40877 37244
rect 40083 37213 40095 37216
rect 40037 37207 40095 37213
rect 40865 37213 40877 37216
rect 40911 37244 40923 37247
rect 40954 37244 40960 37256
rect 40911 37216 40960 37244
rect 40911 37213 40923 37216
rect 40865 37207 40923 37213
rect 40954 37204 40960 37216
rect 41012 37204 41018 37256
rect 41693 37247 41751 37253
rect 41693 37244 41705 37247
rect 41386 37216 41705 37244
rect 28718 37176 28724 37188
rect 28679 37148 28724 37176
rect 28718 37136 28724 37148
rect 28776 37136 28782 37188
rect 30926 37136 30932 37188
rect 30984 37176 30990 37188
rect 31846 37176 31852 37188
rect 30984 37148 31852 37176
rect 30984 37136 30990 37148
rect 31846 37136 31852 37148
rect 31904 37136 31910 37188
rect 40221 37179 40279 37185
rect 40221 37145 40233 37179
rect 40267 37176 40279 37179
rect 41386 37176 41414 37216
rect 41693 37213 41705 37216
rect 41739 37213 41751 37247
rect 43990 37244 43996 37256
rect 43951 37216 43996 37244
rect 41693 37207 41751 37213
rect 43990 37204 43996 37216
rect 44048 37204 44054 37256
rect 44100 37253 44128 37340
rect 44085 37247 44143 37253
rect 44085 37213 44097 37247
rect 44131 37213 44143 37247
rect 44266 37244 44272 37256
rect 44227 37216 44272 37244
rect 44085 37207 44143 37213
rect 40267 37148 41414 37176
rect 40267 37145 40279 37148
rect 40221 37139 40279 37145
rect 43806 37136 43812 37188
rect 43864 37176 43870 37188
rect 44100 37176 44128 37207
rect 44266 37204 44272 37216
rect 44324 37204 44330 37256
rect 46290 37244 46296 37256
rect 46251 37216 46296 37244
rect 46290 37204 46296 37216
rect 46348 37204 46354 37256
rect 43864 37148 44128 37176
rect 46477 37179 46535 37185
rect 43864 37136 43870 37148
rect 46477 37145 46489 37179
rect 46523 37176 46535 37179
rect 47486 37176 47492 37188
rect 46523 37148 47492 37176
rect 46523 37145 46535 37148
rect 46477 37139 46535 37145
rect 47486 37136 47492 37148
rect 47544 37136 47550 37188
rect 48130 37176 48136 37188
rect 48091 37148 48136 37176
rect 48130 37136 48136 37148
rect 48188 37136 48194 37188
rect 24670 37068 24676 37120
rect 24728 37108 24734 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24728 37080 24777 37108
rect 24728 37068 24734 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 27246 37068 27252 37120
rect 27304 37108 27310 37120
rect 27617 37111 27675 37117
rect 27617 37108 27629 37111
rect 27304 37080 27629 37108
rect 27304 37068 27310 37080
rect 27617 37077 27629 37080
rect 27663 37077 27675 37111
rect 28350 37108 28356 37120
rect 28311 37080 28356 37108
rect 27617 37071 27675 37077
rect 28350 37068 28356 37080
rect 28408 37068 28414 37120
rect 35069 37111 35127 37117
rect 35069 37077 35081 37111
rect 35115 37108 35127 37111
rect 35434 37108 35440 37120
rect 35115 37080 35440 37108
rect 35115 37077 35127 37080
rect 35069 37071 35127 37077
rect 35434 37068 35440 37080
rect 35492 37068 35498 37120
rect 35989 37111 36047 37117
rect 35989 37077 36001 37111
rect 36035 37108 36047 37111
rect 36354 37108 36360 37120
rect 36035 37080 36360 37108
rect 36035 37077 36047 37080
rect 35989 37071 36047 37077
rect 36354 37068 36360 37080
rect 36412 37068 36418 37120
rect 36906 37108 36912 37120
rect 36867 37080 36912 37108
rect 36906 37068 36912 37080
rect 36964 37068 36970 37120
rect 41049 37111 41107 37117
rect 41049 37077 41061 37111
rect 41095 37108 41107 37111
rect 41414 37108 41420 37120
rect 41095 37080 41420 37108
rect 41095 37077 41107 37080
rect 41049 37071 41107 37077
rect 41414 37068 41420 37080
rect 41472 37068 41478 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 36173 36907 36231 36913
rect 36173 36873 36185 36907
rect 36219 36904 36231 36907
rect 36906 36904 36912 36916
rect 36219 36876 36912 36904
rect 36219 36873 36231 36876
rect 36173 36867 36231 36873
rect 36906 36864 36912 36876
rect 36964 36864 36970 36916
rect 27614 36836 27620 36848
rect 26988 36808 27620 36836
rect 24302 36777 24308 36780
rect 24296 36731 24308 36777
rect 24360 36768 24366 36780
rect 26988 36777 27016 36808
rect 27614 36796 27620 36808
rect 27672 36836 27678 36848
rect 27890 36836 27896 36848
rect 27672 36808 27896 36836
rect 27672 36796 27678 36808
rect 27890 36796 27896 36808
rect 27948 36796 27954 36848
rect 28350 36796 28356 36848
rect 28408 36836 28414 36848
rect 29058 36839 29116 36845
rect 29058 36836 29070 36839
rect 28408 36808 29070 36836
rect 28408 36796 28414 36808
rect 29058 36805 29070 36808
rect 29104 36805 29116 36839
rect 44726 36836 44732 36848
rect 29058 36799 29116 36805
rect 34256 36808 35388 36836
rect 44687 36808 44732 36836
rect 27246 36777 27252 36780
rect 26973 36771 27031 36777
rect 24360 36740 24396 36768
rect 24302 36728 24308 36731
rect 24360 36728 24366 36740
rect 26973 36737 26985 36771
rect 27019 36737 27031 36771
rect 27240 36768 27252 36777
rect 27207 36740 27252 36768
rect 26973 36731 27031 36737
rect 27240 36731 27252 36740
rect 27246 36728 27252 36731
rect 27304 36728 27310 36780
rect 27908 36768 27936 36796
rect 33134 36777 33140 36780
rect 28813 36771 28871 36777
rect 28813 36768 28825 36771
rect 27908 36740 28825 36768
rect 28813 36737 28825 36740
rect 28859 36737 28871 36771
rect 28813 36731 28871 36737
rect 33128 36731 33140 36777
rect 33192 36768 33198 36780
rect 33192 36740 33228 36768
rect 33134 36728 33140 36731
rect 33192 36728 33198 36740
rect 24029 36703 24087 36709
rect 24029 36669 24041 36703
rect 24075 36669 24087 36703
rect 24029 36663 24087 36669
rect 24044 36564 24072 36663
rect 31754 36660 31760 36712
rect 31812 36700 31818 36712
rect 32122 36700 32128 36712
rect 31812 36672 32128 36700
rect 31812 36660 31818 36672
rect 32122 36660 32128 36672
rect 32180 36700 32186 36712
rect 32861 36703 32919 36709
rect 32861 36700 32873 36703
rect 32180 36672 32873 36700
rect 32180 36660 32186 36672
rect 32861 36669 32873 36672
rect 32907 36669 32919 36703
rect 32861 36663 32919 36669
rect 34256 36576 34284 36808
rect 35360 36777 35388 36808
rect 44726 36796 44732 36808
rect 44784 36796 44790 36848
rect 44945 36839 45003 36845
rect 44945 36805 44957 36839
rect 44991 36836 45003 36839
rect 46198 36836 46204 36848
rect 44991 36808 46204 36836
rect 44991 36805 45003 36808
rect 44945 36799 45003 36805
rect 46198 36796 46204 36808
rect 46256 36796 46262 36848
rect 46290 36796 46296 36848
rect 46348 36836 46354 36848
rect 46348 36808 47808 36836
rect 46348 36796 46354 36808
rect 34977 36771 35035 36777
rect 34977 36737 34989 36771
rect 35023 36737 35035 36771
rect 34977 36731 35035 36737
rect 35069 36771 35127 36777
rect 35069 36737 35081 36771
rect 35115 36737 35127 36771
rect 35069 36731 35127 36737
rect 35253 36771 35311 36777
rect 35253 36737 35265 36771
rect 35299 36737 35311 36771
rect 35253 36731 35311 36737
rect 35345 36771 35403 36777
rect 35345 36737 35357 36771
rect 35391 36737 35403 36771
rect 35986 36768 35992 36780
rect 35947 36740 35992 36768
rect 35345 36731 35403 36737
rect 24394 36564 24400 36576
rect 24044 36536 24400 36564
rect 24394 36524 24400 36536
rect 24452 36564 24458 36576
rect 24762 36564 24768 36576
rect 24452 36536 24768 36564
rect 24452 36524 24458 36536
rect 24762 36524 24768 36536
rect 24820 36524 24826 36576
rect 25406 36564 25412 36576
rect 25367 36536 25412 36564
rect 25406 36524 25412 36536
rect 25464 36524 25470 36576
rect 27154 36524 27160 36576
rect 27212 36564 27218 36576
rect 28353 36567 28411 36573
rect 28353 36564 28365 36567
rect 27212 36536 28365 36564
rect 27212 36524 27218 36536
rect 28353 36533 28365 36536
rect 28399 36533 28411 36567
rect 30190 36564 30196 36576
rect 30151 36536 30196 36564
rect 28353 36527 28411 36533
rect 30190 36524 30196 36536
rect 30248 36524 30254 36576
rect 34238 36564 34244 36576
rect 34199 36536 34244 36564
rect 34238 36524 34244 36536
rect 34296 36524 34302 36576
rect 34514 36524 34520 36576
rect 34572 36564 34578 36576
rect 34793 36567 34851 36573
rect 34793 36564 34805 36567
rect 34572 36536 34805 36564
rect 34572 36524 34578 36536
rect 34793 36533 34805 36536
rect 34839 36533 34851 36567
rect 34992 36564 35020 36731
rect 35084 36632 35112 36731
rect 35268 36700 35296 36731
rect 35986 36728 35992 36740
rect 36044 36728 36050 36780
rect 36262 36768 36268 36780
rect 36223 36740 36268 36768
rect 36262 36728 36268 36740
rect 36320 36728 36326 36780
rect 39025 36771 39083 36777
rect 39025 36737 39037 36771
rect 39071 36768 39083 36771
rect 39850 36768 39856 36780
rect 39071 36740 39856 36768
rect 39071 36737 39083 36740
rect 39025 36731 39083 36737
rect 39850 36728 39856 36740
rect 39908 36728 39914 36780
rect 41414 36728 41420 36780
rect 41472 36768 41478 36780
rect 47026 36768 47032 36780
rect 41472 36740 41517 36768
rect 46987 36740 47032 36768
rect 41472 36728 41478 36740
rect 47026 36728 47032 36740
rect 47084 36728 47090 36780
rect 47780 36777 47808 36808
rect 47765 36771 47823 36777
rect 47765 36737 47777 36771
rect 47811 36737 47823 36771
rect 47765 36731 47823 36737
rect 36004 36700 36032 36728
rect 35268 36672 36032 36700
rect 35618 36632 35624 36644
rect 35084 36604 35624 36632
rect 35618 36592 35624 36604
rect 35676 36592 35682 36644
rect 36262 36632 36268 36644
rect 35728 36604 36268 36632
rect 35342 36564 35348 36576
rect 34992 36536 35348 36564
rect 34793 36527 34851 36533
rect 35342 36524 35348 36536
rect 35400 36564 35406 36576
rect 35728 36564 35756 36604
rect 36262 36592 36268 36604
rect 36320 36592 36326 36644
rect 40402 36592 40408 36644
rect 40460 36632 40466 36644
rect 43990 36632 43996 36644
rect 40460 36604 43996 36632
rect 40460 36592 40466 36604
rect 43990 36592 43996 36604
rect 44048 36592 44054 36644
rect 44174 36592 44180 36644
rect 44232 36632 44238 36644
rect 45097 36635 45155 36641
rect 45097 36632 45109 36635
rect 44232 36604 45109 36632
rect 44232 36592 44238 36604
rect 45097 36601 45109 36604
rect 45143 36601 45155 36635
rect 45097 36595 45155 36601
rect 35400 36536 35756 36564
rect 35400 36524 35406 36536
rect 35802 36524 35808 36576
rect 35860 36564 35866 36576
rect 40494 36564 40500 36576
rect 35860 36536 35905 36564
rect 40455 36536 40500 36564
rect 35860 36524 35866 36536
rect 40494 36524 40500 36536
rect 40552 36524 40558 36576
rect 41230 36564 41236 36576
rect 41191 36536 41236 36564
rect 41230 36524 41236 36536
rect 41288 36524 41294 36576
rect 44913 36567 44971 36573
rect 44913 36533 44925 36567
rect 44959 36564 44971 36567
rect 45186 36564 45192 36576
rect 44959 36536 45192 36564
rect 44959 36533 44971 36536
rect 44913 36527 44971 36533
rect 45186 36524 45192 36536
rect 45244 36524 45250 36576
rect 45830 36524 45836 36576
rect 45888 36564 45894 36576
rect 46658 36564 46664 36576
rect 45888 36536 46664 36564
rect 45888 36524 45894 36536
rect 46658 36524 46664 36536
rect 46716 36524 46722 36576
rect 46842 36564 46848 36576
rect 46803 36536 46848 36564
rect 46842 36524 46848 36536
rect 46900 36524 46906 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 25774 36360 25780 36372
rect 25735 36332 25780 36360
rect 25774 36320 25780 36332
rect 25832 36360 25838 36372
rect 25832 36332 26234 36360
rect 25832 36320 25838 36332
rect 26206 36292 26234 36332
rect 26878 36320 26884 36372
rect 26936 36360 26942 36372
rect 42242 36360 42248 36372
rect 26936 36332 42104 36360
rect 42203 36332 42248 36360
rect 26936 36320 26942 36332
rect 26789 36295 26847 36301
rect 26789 36292 26801 36295
rect 26206 36264 26801 36292
rect 26789 36261 26801 36264
rect 26835 36292 26847 36295
rect 27246 36292 27252 36304
rect 26835 36264 27252 36292
rect 26835 36261 26847 36264
rect 26789 36255 26847 36261
rect 27246 36252 27252 36264
rect 27304 36252 27310 36304
rect 40402 36292 40408 36304
rect 40363 36264 40408 36292
rect 40402 36252 40408 36264
rect 40460 36252 40466 36304
rect 42076 36292 42104 36332
rect 42242 36320 42248 36332
rect 42300 36320 42306 36372
rect 45830 36360 45836 36372
rect 42352 36332 45836 36360
rect 42352 36292 42380 36332
rect 45830 36320 45836 36332
rect 45888 36320 45894 36372
rect 46198 36320 46204 36372
rect 46256 36360 46262 36372
rect 46293 36363 46351 36369
rect 46293 36360 46305 36363
rect 46256 36332 46305 36360
rect 46256 36320 46262 36332
rect 46293 36329 46305 36332
rect 46339 36329 46351 36363
rect 46934 36360 46940 36372
rect 46293 36323 46351 36329
rect 46768 36332 46940 36360
rect 42076 36264 42380 36292
rect 45741 36295 45799 36301
rect 45741 36261 45753 36295
rect 45787 36292 45799 36295
rect 46768 36292 46796 36332
rect 46934 36320 46940 36332
rect 46992 36320 46998 36372
rect 45787 36264 46796 36292
rect 45787 36261 45799 36264
rect 45741 36255 45799 36261
rect 29178 36184 29184 36236
rect 29236 36224 29242 36236
rect 29549 36227 29607 36233
rect 29549 36224 29561 36227
rect 29236 36196 29561 36224
rect 29236 36184 29242 36196
rect 29549 36193 29561 36196
rect 29595 36224 29607 36227
rect 30190 36224 30196 36236
rect 29595 36196 30196 36224
rect 29595 36193 29607 36196
rect 29549 36187 29607 36193
rect 30190 36184 30196 36196
rect 30248 36184 30254 36236
rect 34238 36184 34244 36236
rect 34296 36224 34302 36236
rect 34701 36227 34759 36233
rect 34701 36224 34713 36227
rect 34296 36196 34713 36224
rect 34296 36184 34302 36196
rect 34701 36193 34713 36196
rect 34747 36193 34759 36227
rect 36446 36224 36452 36236
rect 36407 36196 36452 36224
rect 34701 36187 34759 36193
rect 36446 36184 36452 36196
rect 36504 36184 36510 36236
rect 45554 36184 45560 36236
rect 45612 36224 45618 36236
rect 46750 36224 46756 36236
rect 45612 36196 46756 36224
rect 45612 36184 45618 36196
rect 46750 36184 46756 36196
rect 46808 36184 46814 36236
rect 19889 36159 19947 36165
rect 19889 36125 19901 36159
rect 19935 36156 19947 36159
rect 19978 36156 19984 36168
rect 19935 36128 19984 36156
rect 19935 36125 19947 36128
rect 19889 36119 19947 36125
rect 19978 36116 19984 36128
rect 20036 36156 20042 36168
rect 24394 36156 24400 36168
rect 20036 36128 22048 36156
rect 24355 36128 24400 36156
rect 20036 36116 20042 36128
rect 20349 36091 20407 36097
rect 20349 36057 20361 36091
rect 20395 36057 20407 36091
rect 22020 36088 22048 36128
rect 24394 36116 24400 36128
rect 24452 36116 24458 36168
rect 24670 36165 24676 36168
rect 24664 36156 24676 36165
rect 24631 36128 24676 36156
rect 24664 36119 24676 36128
rect 24670 36116 24676 36119
rect 24728 36116 24734 36168
rect 26786 36116 26792 36168
rect 26844 36156 26850 36168
rect 26973 36159 27031 36165
rect 26973 36156 26985 36159
rect 26844 36128 26985 36156
rect 26844 36116 26850 36128
rect 26973 36125 26985 36128
rect 27019 36125 27031 36159
rect 26973 36119 27031 36125
rect 27065 36159 27123 36165
rect 27065 36125 27077 36159
rect 27111 36156 27123 36159
rect 27154 36156 27160 36168
rect 27111 36128 27160 36156
rect 27111 36125 27123 36128
rect 27065 36119 27123 36125
rect 27154 36116 27160 36128
rect 27212 36116 27218 36168
rect 27338 36116 27344 36168
rect 27396 36116 27402 36168
rect 29733 36159 29791 36165
rect 29733 36125 29745 36159
rect 29779 36156 29791 36159
rect 30926 36156 30932 36168
rect 29779 36128 30932 36156
rect 29779 36125 29791 36128
rect 29733 36119 29791 36125
rect 30926 36116 30932 36128
rect 30984 36116 30990 36168
rect 34974 36156 34980 36168
rect 34935 36128 34980 36156
rect 34974 36116 34980 36128
rect 35032 36116 35038 36168
rect 35434 36116 35440 36168
rect 35492 36156 35498 36168
rect 36173 36159 36231 36165
rect 36173 36156 36185 36159
rect 35492 36128 36185 36156
rect 35492 36116 35498 36128
rect 36173 36125 36185 36128
rect 36219 36125 36231 36159
rect 36173 36119 36231 36125
rect 36262 36116 36268 36168
rect 36320 36156 36326 36168
rect 36541 36159 36599 36165
rect 36320 36128 36365 36156
rect 36320 36116 36326 36128
rect 36541 36125 36553 36159
rect 36587 36156 36599 36159
rect 36906 36156 36912 36168
rect 36587 36128 36912 36156
rect 36587 36125 36599 36128
rect 36541 36119 36599 36125
rect 26694 36088 26700 36100
rect 22020 36060 26700 36088
rect 20349 36051 20407 36057
rect 20364 36020 20392 36051
rect 26694 36048 26700 36060
rect 26752 36048 26758 36100
rect 27356 36088 27384 36116
rect 27172 36060 27384 36088
rect 20438 36020 20444 36032
rect 20351 35992 20444 36020
rect 20438 35980 20444 35992
rect 20496 36020 20502 36032
rect 26878 36020 26884 36032
rect 20496 35992 26884 36020
rect 20496 35980 20502 35992
rect 26878 35980 26884 35992
rect 26936 35980 26942 36032
rect 27172 36029 27200 36060
rect 35618 36048 35624 36100
rect 35676 36088 35682 36100
rect 36556 36088 36584 36119
rect 36906 36116 36912 36128
rect 36964 36116 36970 36168
rect 40865 36159 40923 36165
rect 40865 36125 40877 36159
rect 40911 36156 40923 36159
rect 42705 36159 42763 36165
rect 42705 36156 42717 36159
rect 40911 36128 42717 36156
rect 40911 36125 40923 36128
rect 40865 36119 40923 36125
rect 42705 36125 42717 36128
rect 42751 36156 42763 36159
rect 42794 36156 42800 36168
rect 42751 36128 42800 36156
rect 42751 36125 42763 36128
rect 42705 36119 42763 36125
rect 42794 36116 42800 36128
rect 42852 36116 42858 36168
rect 45922 36156 45928 36168
rect 45883 36128 45928 36156
rect 45922 36116 45928 36128
rect 45980 36116 45986 36168
rect 46842 36116 46848 36168
rect 46900 36156 46906 36168
rect 47009 36159 47067 36165
rect 47009 36156 47021 36159
rect 46900 36128 47021 36156
rect 46900 36116 46906 36128
rect 47009 36125 47021 36128
rect 47055 36125 47067 36159
rect 47009 36119 47067 36125
rect 35676 36060 36584 36088
rect 40221 36091 40279 36097
rect 35676 36048 35682 36060
rect 40221 36057 40233 36091
rect 40267 36088 40279 36091
rect 40954 36088 40960 36100
rect 40267 36060 40960 36088
rect 40267 36057 40279 36060
rect 40221 36051 40279 36057
rect 40954 36048 40960 36060
rect 41012 36048 41018 36100
rect 41132 36091 41190 36097
rect 41132 36057 41144 36091
rect 41178 36088 41190 36091
rect 41230 36088 41236 36100
rect 41178 36060 41236 36088
rect 41178 36057 41190 36060
rect 41132 36051 41190 36057
rect 41230 36048 41236 36060
rect 41288 36048 41294 36100
rect 42978 36097 42984 36100
rect 42972 36051 42984 36097
rect 43036 36088 43042 36100
rect 46017 36091 46075 36097
rect 43036 36060 43072 36088
rect 42978 36048 42984 36051
rect 43036 36048 43042 36060
rect 46017 36057 46029 36091
rect 46063 36088 46075 36091
rect 46566 36088 46572 36100
rect 46063 36060 46572 36088
rect 46063 36057 46075 36060
rect 46017 36051 46075 36057
rect 46566 36048 46572 36060
rect 46624 36048 46630 36100
rect 27157 36023 27215 36029
rect 27157 35989 27169 36023
rect 27203 35989 27215 36023
rect 27157 35983 27215 35989
rect 27341 36023 27399 36029
rect 27341 35989 27353 36023
rect 27387 36020 27399 36023
rect 27798 36020 27804 36032
rect 27387 35992 27804 36020
rect 27387 35989 27399 35992
rect 27341 35983 27399 35989
rect 27798 35980 27804 35992
rect 27856 35980 27862 36032
rect 29546 35980 29552 36032
rect 29604 36020 29610 36032
rect 29917 36023 29975 36029
rect 29917 36020 29929 36023
rect 29604 35992 29929 36020
rect 29604 35980 29610 35992
rect 29917 35989 29929 35992
rect 29963 35989 29975 36023
rect 35986 36020 35992 36032
rect 35947 35992 35992 36020
rect 29917 35983 29975 35989
rect 35986 35980 35992 35992
rect 36044 35980 36050 36032
rect 44082 36020 44088 36032
rect 44043 35992 44088 36020
rect 44082 35980 44088 35992
rect 44140 35980 44146 36032
rect 46109 36023 46167 36029
rect 46109 35989 46121 36023
rect 46155 36020 46167 36023
rect 46382 36020 46388 36032
rect 46155 35992 46388 36020
rect 46155 35989 46167 35992
rect 46109 35983 46167 35989
rect 46382 35980 46388 35992
rect 46440 36020 46446 36032
rect 48133 36023 48191 36029
rect 48133 36020 48145 36023
rect 46440 35992 48145 36020
rect 46440 35980 46446 35992
rect 48133 35989 48145 35992
rect 48179 35989 48191 36023
rect 48133 35983 48191 35989
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 24213 35819 24271 35825
rect 24213 35785 24225 35819
rect 24259 35816 24271 35819
rect 24302 35816 24308 35828
rect 24259 35788 24308 35816
rect 24259 35785 24271 35788
rect 24213 35779 24271 35785
rect 24302 35776 24308 35788
rect 24360 35776 24366 35828
rect 24946 35776 24952 35828
rect 25004 35816 25010 35828
rect 25225 35819 25283 35825
rect 25225 35816 25237 35819
rect 25004 35788 25237 35816
rect 25004 35776 25010 35788
rect 25225 35785 25237 35788
rect 25271 35785 25283 35819
rect 25225 35779 25283 35785
rect 36998 35776 37004 35828
rect 37056 35816 37062 35828
rect 39853 35819 39911 35825
rect 39853 35816 39865 35819
rect 37056 35788 39865 35816
rect 37056 35776 37062 35788
rect 39853 35785 39865 35788
rect 39899 35785 39911 35819
rect 40678 35816 40684 35828
rect 40639 35788 40684 35816
rect 39853 35779 39911 35785
rect 40678 35776 40684 35788
rect 40736 35776 40742 35828
rect 42797 35819 42855 35825
rect 42797 35785 42809 35819
rect 42843 35816 42855 35819
rect 42978 35816 42984 35828
rect 42843 35788 42984 35816
rect 42843 35785 42855 35788
rect 42797 35779 42855 35785
rect 42978 35776 42984 35788
rect 43036 35776 43042 35828
rect 43901 35819 43959 35825
rect 43901 35785 43913 35819
rect 43947 35816 43959 35819
rect 44082 35816 44088 35828
rect 43947 35788 44088 35816
rect 43947 35785 43959 35788
rect 43901 35779 43959 35785
rect 44082 35776 44088 35788
rect 44140 35816 44146 35828
rect 46845 35819 46903 35825
rect 46845 35816 46857 35819
rect 44140 35788 45508 35816
rect 44140 35776 44146 35788
rect 25685 35751 25743 35757
rect 25685 35717 25697 35751
rect 25731 35748 25743 35751
rect 26050 35748 26056 35760
rect 25731 35720 26056 35748
rect 25731 35717 25743 35720
rect 25685 35711 25743 35717
rect 26050 35708 26056 35720
rect 26108 35708 26114 35760
rect 26973 35751 27031 35757
rect 26973 35717 26985 35751
rect 27019 35748 27031 35751
rect 27062 35748 27068 35760
rect 27019 35720 27068 35748
rect 27019 35717 27031 35720
rect 26973 35711 27031 35717
rect 27062 35708 27068 35720
rect 27120 35708 27126 35760
rect 36446 35748 36452 35760
rect 35360 35720 36452 35748
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35680 24455 35683
rect 24946 35680 24952 35692
rect 24443 35652 24952 35680
rect 24443 35649 24455 35652
rect 24397 35643 24455 35649
rect 24946 35640 24952 35652
rect 25004 35640 25010 35692
rect 25038 35640 25044 35692
rect 25096 35680 25102 35692
rect 25096 35652 25141 35680
rect 25096 35640 25102 35652
rect 25866 35640 25872 35692
rect 25924 35680 25930 35692
rect 25961 35683 26019 35689
rect 25961 35680 25973 35683
rect 25924 35652 25973 35680
rect 25924 35640 25930 35652
rect 25961 35649 25973 35652
rect 26007 35649 26019 35683
rect 27246 35680 27252 35692
rect 27207 35652 27252 35680
rect 25961 35643 26019 35649
rect 27246 35640 27252 35652
rect 27304 35640 27310 35692
rect 29546 35680 29552 35692
rect 29507 35652 29552 35680
rect 29546 35640 29552 35652
rect 29604 35640 29610 35692
rect 32306 35680 32312 35692
rect 32267 35652 32312 35680
rect 32306 35640 32312 35652
rect 32364 35640 32370 35692
rect 33502 35640 33508 35692
rect 33560 35680 33566 35692
rect 34974 35680 34980 35692
rect 33560 35652 34980 35680
rect 33560 35640 33566 35652
rect 34974 35640 34980 35652
rect 35032 35680 35038 35692
rect 35069 35683 35127 35689
rect 35069 35680 35081 35683
rect 35032 35652 35081 35680
rect 35032 35640 35038 35652
rect 35069 35649 35081 35652
rect 35115 35649 35127 35683
rect 35250 35680 35256 35692
rect 35211 35652 35256 35680
rect 35069 35643 35127 35649
rect 35250 35640 35256 35652
rect 35308 35640 35314 35692
rect 35360 35689 35388 35720
rect 36446 35708 36452 35720
rect 36504 35708 36510 35760
rect 39209 35751 39267 35757
rect 39209 35717 39221 35751
rect 39255 35748 39267 35751
rect 39669 35751 39727 35757
rect 39669 35748 39681 35751
rect 39255 35720 39681 35748
rect 39255 35717 39267 35720
rect 39209 35711 39267 35717
rect 39669 35717 39681 35720
rect 39715 35717 39727 35751
rect 43990 35748 43996 35760
rect 43903 35720 43996 35748
rect 39669 35711 39727 35717
rect 43990 35708 43996 35720
rect 44048 35748 44054 35760
rect 44358 35748 44364 35760
rect 44048 35720 44364 35748
rect 44048 35708 44054 35720
rect 44358 35708 44364 35720
rect 44416 35708 44422 35760
rect 45480 35757 45508 35788
rect 45572 35788 46857 35816
rect 45465 35751 45523 35757
rect 45465 35717 45477 35751
rect 45511 35717 45523 35751
rect 45465 35711 45523 35717
rect 35345 35683 35403 35689
rect 35345 35649 35357 35683
rect 35391 35649 35403 35683
rect 35345 35643 35403 35649
rect 35434 35640 35440 35692
rect 35492 35680 35498 35692
rect 35492 35652 35537 35680
rect 35492 35640 35498 35652
rect 35618 35640 35624 35692
rect 35676 35680 35682 35692
rect 38930 35680 38936 35692
rect 35676 35652 35721 35680
rect 38891 35652 38936 35680
rect 35676 35640 35682 35652
rect 38930 35640 38936 35652
rect 38988 35640 38994 35692
rect 39942 35640 39948 35692
rect 40000 35680 40006 35692
rect 40862 35680 40868 35692
rect 40000 35652 40045 35680
rect 40823 35652 40868 35680
rect 40000 35640 40006 35652
rect 40862 35640 40868 35652
rect 40920 35640 40926 35692
rect 42978 35680 42984 35692
rect 42939 35652 42984 35680
rect 42978 35640 42984 35652
rect 43036 35640 43042 35692
rect 43625 35683 43683 35689
rect 43625 35649 43637 35683
rect 43671 35680 43683 35683
rect 44545 35683 44603 35689
rect 44545 35680 44557 35683
rect 43671 35652 44557 35680
rect 43671 35649 43683 35652
rect 43625 35643 43683 35649
rect 44545 35649 44557 35652
rect 44591 35649 44603 35683
rect 44545 35643 44603 35649
rect 44634 35640 44640 35692
rect 44692 35680 44698 35692
rect 44729 35683 44787 35689
rect 44729 35680 44741 35683
rect 44692 35652 44741 35680
rect 44692 35640 44698 35652
rect 44729 35649 44741 35652
rect 44775 35649 44787 35683
rect 44729 35643 44787 35649
rect 44913 35683 44971 35689
rect 44913 35649 44925 35683
rect 44959 35680 44971 35683
rect 44959 35678 45416 35680
rect 45572 35678 45600 35788
rect 46845 35785 46857 35788
rect 46891 35785 46903 35819
rect 46845 35779 46903 35785
rect 47026 35776 47032 35828
rect 47084 35816 47090 35828
rect 47949 35819 48007 35825
rect 47949 35816 47961 35819
rect 47084 35788 47961 35816
rect 47084 35776 47090 35788
rect 47949 35785 47961 35788
rect 47995 35785 48007 35819
rect 47949 35779 48007 35785
rect 45738 35680 45744 35692
rect 44959 35652 45600 35678
rect 45699 35652 45744 35680
rect 44959 35649 44971 35652
rect 45388 35650 45600 35652
rect 44913 35643 44971 35649
rect 45738 35640 45744 35652
rect 45796 35640 45802 35692
rect 46382 35680 46388 35692
rect 46343 35652 46388 35680
rect 46382 35640 46388 35652
rect 46440 35640 46446 35692
rect 46661 35683 46719 35689
rect 46661 35649 46673 35683
rect 46707 35680 46719 35683
rect 46934 35680 46940 35692
rect 46707 35652 46940 35680
rect 46707 35649 46719 35652
rect 46661 35643 46719 35649
rect 46934 35640 46940 35652
rect 46992 35680 46998 35692
rect 47581 35683 47639 35689
rect 47581 35680 47593 35683
rect 46992 35652 47593 35680
rect 46992 35640 46998 35652
rect 47581 35649 47593 35652
rect 47627 35649 47639 35683
rect 47762 35680 47768 35692
rect 47723 35652 47768 35680
rect 47581 35643 47639 35649
rect 47762 35640 47768 35652
rect 47820 35640 47826 35692
rect 24857 35615 24915 35621
rect 24857 35581 24869 35615
rect 24903 35612 24915 35615
rect 25406 35612 25412 35624
rect 24903 35584 25412 35612
rect 24903 35581 24915 35584
rect 24857 35575 24915 35581
rect 25406 35572 25412 35584
rect 25464 35572 25470 35624
rect 25498 35572 25504 35624
rect 25556 35612 25562 35624
rect 25777 35615 25835 35621
rect 25777 35612 25789 35615
rect 25556 35584 25789 35612
rect 25556 35572 25562 35584
rect 25777 35581 25789 35584
rect 25823 35581 25835 35615
rect 27154 35612 27160 35624
rect 27115 35584 27160 35612
rect 25777 35575 25835 35581
rect 27154 35572 27160 35584
rect 27212 35572 27218 35624
rect 32401 35615 32459 35621
rect 32401 35581 32413 35615
rect 32447 35612 32459 35615
rect 33226 35612 33232 35624
rect 32447 35584 33232 35612
rect 32447 35581 32459 35584
rect 32401 35575 32459 35581
rect 33226 35572 33232 35584
rect 33284 35572 33290 35624
rect 38562 35572 38568 35624
rect 38620 35612 38626 35624
rect 39209 35615 39267 35621
rect 39209 35612 39221 35615
rect 38620 35584 39221 35612
rect 38620 35572 38626 35584
rect 39209 35581 39221 35584
rect 39255 35581 39267 35615
rect 43714 35612 43720 35624
rect 43675 35584 43720 35612
rect 39209 35575 39267 35581
rect 43714 35572 43720 35584
rect 43772 35572 43778 35624
rect 44085 35615 44143 35621
rect 44085 35581 44097 35615
rect 44131 35612 44143 35615
rect 44174 35612 44180 35624
rect 44131 35584 44180 35612
rect 44131 35581 44143 35584
rect 44085 35575 44143 35581
rect 44174 35572 44180 35584
rect 44232 35572 44238 35624
rect 45005 35615 45063 35621
rect 45005 35581 45017 35615
rect 45051 35581 45063 35615
rect 45005 35575 45063 35581
rect 25424 35544 25452 35572
rect 26786 35544 26792 35556
rect 25424 35516 26792 35544
rect 26786 35504 26792 35516
rect 26844 35544 26850 35556
rect 26844 35516 27016 35544
rect 26844 35504 26850 35516
rect 25682 35436 25688 35488
rect 25740 35476 25746 35488
rect 25958 35476 25964 35488
rect 25740 35448 25964 35476
rect 25740 35436 25746 35448
rect 25958 35436 25964 35448
rect 26016 35436 26022 35488
rect 26142 35476 26148 35488
rect 26103 35448 26148 35476
rect 26142 35436 26148 35448
rect 26200 35436 26206 35488
rect 26988 35485 27016 35516
rect 28718 35504 28724 35556
rect 28776 35544 28782 35556
rect 32122 35544 32128 35556
rect 28776 35516 32128 35544
rect 28776 35504 28782 35516
rect 32122 35504 32128 35516
rect 32180 35544 32186 35556
rect 40402 35544 40408 35556
rect 32180 35516 40408 35544
rect 32180 35504 32186 35516
rect 40402 35504 40408 35516
rect 40460 35504 40466 35556
rect 45020 35544 45048 35575
rect 45186 35572 45192 35624
rect 45244 35612 45250 35624
rect 45557 35615 45615 35621
rect 45557 35612 45569 35615
rect 45244 35584 45569 35612
rect 45244 35572 45250 35584
rect 45557 35581 45569 35584
rect 45603 35581 45615 35615
rect 46566 35612 46572 35624
rect 46527 35584 46572 35612
rect 45557 35575 45615 35581
rect 46566 35572 46572 35584
rect 46624 35572 46630 35624
rect 45925 35547 45983 35553
rect 45925 35544 45937 35547
rect 45020 35516 45937 35544
rect 45925 35513 45937 35516
rect 45971 35513 45983 35547
rect 45925 35507 45983 35513
rect 26973 35479 27031 35485
rect 26973 35445 26985 35479
rect 27019 35445 27031 35479
rect 26973 35439 27031 35445
rect 27062 35436 27068 35488
rect 27120 35476 27126 35488
rect 27433 35479 27491 35485
rect 27433 35476 27445 35479
rect 27120 35448 27445 35476
rect 27120 35436 27126 35448
rect 27433 35445 27445 35448
rect 27479 35445 27491 35479
rect 27433 35439 27491 35445
rect 28994 35436 29000 35488
rect 29052 35476 29058 35488
rect 29362 35476 29368 35488
rect 29052 35448 29368 35476
rect 29052 35436 29058 35448
rect 29362 35436 29368 35448
rect 29420 35436 29426 35488
rect 32214 35436 32220 35488
rect 32272 35476 32278 35488
rect 32677 35479 32735 35485
rect 32677 35476 32689 35479
rect 32272 35448 32689 35476
rect 32272 35436 32278 35448
rect 32677 35445 32689 35448
rect 32723 35445 32735 35479
rect 32677 35439 32735 35445
rect 34698 35436 34704 35488
rect 34756 35476 34762 35488
rect 35805 35479 35863 35485
rect 35805 35476 35817 35479
rect 34756 35448 35817 35476
rect 34756 35436 34762 35448
rect 35805 35445 35817 35448
rect 35851 35445 35863 35479
rect 35805 35439 35863 35445
rect 37366 35436 37372 35488
rect 37424 35476 37430 35488
rect 39025 35479 39083 35485
rect 39025 35476 39037 35479
rect 37424 35448 39037 35476
rect 37424 35436 37430 35448
rect 39025 35445 39037 35448
rect 39071 35445 39083 35479
rect 39025 35439 39083 35445
rect 39669 35479 39727 35485
rect 39669 35445 39681 35479
rect 39715 35476 39727 35479
rect 40126 35476 40132 35488
rect 39715 35448 40132 35476
rect 39715 35445 39727 35448
rect 39669 35439 39727 35445
rect 40126 35436 40132 35448
rect 40184 35436 40190 35488
rect 43438 35476 43444 35488
rect 43399 35448 43444 35476
rect 43438 35436 43444 35448
rect 43496 35436 43502 35488
rect 44726 35436 44732 35488
rect 44784 35476 44790 35488
rect 45465 35479 45523 35485
rect 45465 35476 45477 35479
rect 44784 35448 45477 35476
rect 44784 35436 44790 35448
rect 45465 35445 45477 35448
rect 45511 35445 45523 35479
rect 45465 35439 45523 35445
rect 46014 35436 46020 35488
rect 46072 35476 46078 35488
rect 46385 35479 46443 35485
rect 46385 35476 46397 35479
rect 46072 35448 46397 35476
rect 46072 35436 46078 35448
rect 46385 35445 46397 35448
rect 46431 35445 46443 35479
rect 46385 35439 46443 35445
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 24946 35232 24952 35284
rect 25004 35272 25010 35284
rect 25225 35275 25283 35281
rect 25225 35272 25237 35275
rect 25004 35244 25237 35272
rect 25004 35232 25010 35244
rect 25225 35241 25237 35244
rect 25271 35241 25283 35275
rect 25225 35235 25283 35241
rect 33410 35232 33416 35284
rect 33468 35272 33474 35284
rect 38654 35272 38660 35284
rect 33468 35244 38660 35272
rect 33468 35232 33474 35244
rect 38654 35232 38660 35244
rect 38712 35272 38718 35284
rect 38712 35244 38884 35272
rect 38712 35232 38718 35244
rect 35897 35207 35955 35213
rect 35897 35173 35909 35207
rect 35943 35173 35955 35207
rect 35897 35167 35955 35173
rect 24857 35139 24915 35145
rect 24857 35105 24869 35139
rect 24903 35136 24915 35139
rect 24903 35108 25544 35136
rect 24903 35105 24915 35108
rect 24857 35099 24915 35105
rect 25516 35080 25544 35108
rect 26050 35096 26056 35148
rect 26108 35136 26114 35148
rect 35912 35136 35940 35167
rect 38856 35145 38884 35244
rect 42978 35232 42984 35284
rect 43036 35272 43042 35284
rect 44177 35275 44235 35281
rect 44177 35272 44189 35275
rect 43036 35244 44189 35272
rect 43036 35232 43042 35244
rect 44177 35241 44189 35244
rect 44223 35241 44235 35275
rect 44177 35235 44235 35241
rect 46566 35232 46572 35284
rect 46624 35272 46630 35284
rect 48133 35275 48191 35281
rect 48133 35272 48145 35275
rect 46624 35244 48145 35272
rect 46624 35232 46630 35244
rect 48133 35241 48145 35244
rect 48179 35241 48191 35275
rect 48133 35235 48191 35241
rect 38841 35139 38899 35145
rect 26108 35108 26280 35136
rect 35912 35108 36400 35136
rect 26108 35096 26114 35108
rect 2038 35028 2044 35080
rect 2096 35068 2102 35080
rect 2317 35071 2375 35077
rect 2317 35068 2329 35071
rect 2096 35040 2329 35068
rect 2096 35028 2102 35040
rect 2317 35037 2329 35040
rect 2363 35037 2375 35071
rect 25038 35068 25044 35080
rect 2317 35031 2375 35037
rect 24872 35040 25044 35068
rect 24872 35012 24900 35040
rect 25038 35028 25044 35040
rect 25096 35028 25102 35080
rect 25498 35028 25504 35080
rect 25556 35068 25562 35080
rect 26252 35077 26280 35108
rect 26145 35071 26203 35077
rect 26145 35068 26157 35071
rect 25556 35040 26157 35068
rect 25556 35028 25562 35040
rect 26145 35037 26157 35040
rect 26191 35037 26203 35071
rect 26145 35031 26203 35037
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35037 26295 35071
rect 26237 35031 26295 35037
rect 26421 35071 26479 35077
rect 26421 35037 26433 35071
rect 26467 35068 26479 35071
rect 27709 35071 27767 35077
rect 27709 35068 27721 35071
rect 26467 35040 27721 35068
rect 26467 35037 26479 35040
rect 26421 35031 26479 35037
rect 27709 35037 27721 35040
rect 27755 35037 27767 35071
rect 27709 35031 27767 35037
rect 27798 35028 27804 35080
rect 27856 35068 27862 35080
rect 28169 35071 28227 35077
rect 27856 35040 27901 35068
rect 27856 35028 27862 35040
rect 28169 35037 28181 35071
rect 28215 35068 28227 35071
rect 28994 35068 29000 35080
rect 28215 35040 29000 35068
rect 28215 35037 28227 35040
rect 28169 35031 28227 35037
rect 28994 35028 29000 35040
rect 29052 35028 29058 35080
rect 30929 35071 30987 35077
rect 30929 35037 30941 35071
rect 30975 35068 30987 35071
rect 31754 35068 31760 35080
rect 30975 35040 31760 35068
rect 30975 35037 30987 35040
rect 30929 35031 30987 35037
rect 31754 35028 31760 35040
rect 31812 35028 31818 35080
rect 34698 35068 34704 35080
rect 34659 35040 34704 35068
rect 34698 35028 34704 35040
rect 34756 35028 34762 35080
rect 34882 35068 34888 35080
rect 34843 35040 34888 35068
rect 34882 35028 34888 35040
rect 34940 35028 34946 35080
rect 36170 35068 36176 35080
rect 36131 35040 36176 35068
rect 36170 35028 36176 35040
rect 36228 35028 36234 35080
rect 24854 34960 24860 35012
rect 24912 34960 24918 35012
rect 25866 35000 25872 35012
rect 25827 34972 25872 35000
rect 25866 34960 25872 34972
rect 25924 34960 25930 35012
rect 27893 35003 27951 35009
rect 27893 34969 27905 35003
rect 27939 34969 27951 35003
rect 27893 34963 27951 34969
rect 25958 34892 25964 34944
rect 26016 34932 26022 34944
rect 26053 34935 26111 34941
rect 26053 34932 26065 34935
rect 26016 34904 26065 34932
rect 26016 34892 26022 34904
rect 26053 34901 26065 34904
rect 26099 34901 26111 34935
rect 27522 34932 27528 34944
rect 27483 34904 27528 34932
rect 26053 34895 26111 34901
rect 27522 34892 27528 34904
rect 27580 34892 27586 34944
rect 27908 34932 27936 34963
rect 27982 34960 27988 35012
rect 28040 35009 28046 35012
rect 28040 35003 28069 35009
rect 28057 34969 28069 35003
rect 28040 34963 28069 34969
rect 31196 35003 31254 35009
rect 31196 34969 31208 35003
rect 31242 35000 31254 35003
rect 32858 35000 32864 35012
rect 31242 34972 32864 35000
rect 31242 34969 31254 34972
rect 31196 34963 31254 34969
rect 28040 34960 28046 34963
rect 32858 34960 32864 34972
rect 32916 34960 32922 35012
rect 35894 35000 35900 35012
rect 35855 34972 35900 35000
rect 35894 34960 35900 34972
rect 35952 34960 35958 35012
rect 36372 35000 36400 35108
rect 38841 35105 38853 35139
rect 38887 35105 38899 35139
rect 38841 35099 38899 35105
rect 39114 35096 39120 35148
rect 39172 35136 39178 35148
rect 39301 35139 39359 35145
rect 39301 35136 39313 35139
rect 39172 35108 39313 35136
rect 39172 35096 39178 35108
rect 39301 35105 39313 35108
rect 39347 35105 39359 35139
rect 39301 35099 39359 35105
rect 39408 35108 39896 35136
rect 36633 35071 36691 35077
rect 36633 35037 36645 35071
rect 36679 35068 36691 35071
rect 36679 35040 38884 35068
rect 36679 35037 36691 35040
rect 36633 35031 36691 35037
rect 36878 35003 36936 35009
rect 36878 35000 36890 35003
rect 36372 34972 36890 35000
rect 36878 34969 36890 34972
rect 36924 34969 36936 35003
rect 38856 35000 38884 35040
rect 38930 35028 38936 35080
rect 38988 35068 38994 35080
rect 38988 35040 39033 35068
rect 38988 35028 38994 35040
rect 39408 35000 39436 35108
rect 39868 35077 39896 35108
rect 43714 35096 43720 35148
rect 43772 35136 43778 35148
rect 43809 35139 43867 35145
rect 43809 35136 43821 35139
rect 43772 35108 43821 35136
rect 43772 35096 43778 35108
rect 43809 35105 43821 35108
rect 43855 35136 43867 35139
rect 45738 35136 45744 35148
rect 43855 35108 45744 35136
rect 43855 35105 43867 35108
rect 43809 35099 43867 35105
rect 45738 35096 45744 35108
rect 45796 35096 45802 35148
rect 46750 35136 46756 35148
rect 46711 35108 46756 35136
rect 46750 35096 46756 35108
rect 46808 35096 46814 35148
rect 39853 35071 39911 35077
rect 39853 35037 39865 35071
rect 39899 35068 39911 35071
rect 40494 35068 40500 35080
rect 39899 35040 40500 35068
rect 39899 35037 39911 35040
rect 39853 35031 39911 35037
rect 40494 35028 40500 35040
rect 40552 35028 40558 35080
rect 43993 35071 44051 35077
rect 43993 35037 44005 35071
rect 44039 35068 44051 35071
rect 44174 35068 44180 35080
rect 44039 35040 44180 35068
rect 44039 35037 44051 35040
rect 43993 35031 44051 35037
rect 44174 35028 44180 35040
rect 44232 35028 44238 35080
rect 44726 35028 44732 35080
rect 44784 35068 44790 35080
rect 45005 35071 45063 35077
rect 45005 35068 45017 35071
rect 44784 35040 45017 35068
rect 44784 35028 44790 35040
rect 45005 35037 45017 35040
rect 45051 35037 45063 35071
rect 45005 35031 45063 35037
rect 45189 35071 45247 35077
rect 45189 35037 45201 35071
rect 45235 35037 45247 35071
rect 45189 35031 45247 35037
rect 46293 35071 46351 35077
rect 46293 35037 46305 35071
rect 46339 35068 46351 35071
rect 46842 35068 46848 35080
rect 46339 35040 46848 35068
rect 46339 35037 46351 35040
rect 46293 35031 46351 35037
rect 40126 35009 40132 35012
rect 40120 35000 40132 35009
rect 38856 34972 39436 35000
rect 40087 34972 40132 35000
rect 36878 34963 36936 34969
rect 40120 34963 40132 34972
rect 40126 34960 40132 34963
rect 40184 34960 40190 35012
rect 44192 35000 44220 35028
rect 45204 35000 45232 35031
rect 46842 35028 46848 35040
rect 46900 35028 46906 35080
rect 46998 35003 47056 35009
rect 46998 35000 47010 35003
rect 44192 34972 45232 35000
rect 46124 34972 47010 35000
rect 28718 34932 28724 34944
rect 27908 34904 28724 34932
rect 28718 34892 28724 34904
rect 28776 34892 28782 34944
rect 32306 34932 32312 34944
rect 32219 34904 32312 34932
rect 32306 34892 32312 34904
rect 32364 34932 32370 34944
rect 32674 34932 32680 34944
rect 32364 34904 32680 34932
rect 32364 34892 32370 34904
rect 32674 34892 32680 34904
rect 32732 34892 32738 34944
rect 34793 34935 34851 34941
rect 34793 34901 34805 34935
rect 34839 34932 34851 34935
rect 34974 34932 34980 34944
rect 34839 34904 34980 34932
rect 34839 34901 34851 34904
rect 34793 34895 34851 34901
rect 34974 34892 34980 34904
rect 35032 34892 35038 34944
rect 35434 34892 35440 34944
rect 35492 34932 35498 34944
rect 36081 34935 36139 34941
rect 36081 34932 36093 34935
rect 35492 34904 36093 34932
rect 35492 34892 35498 34904
rect 36081 34901 36093 34904
rect 36127 34932 36139 34935
rect 36998 34932 37004 34944
rect 36127 34904 37004 34932
rect 36127 34901 36139 34904
rect 36081 34895 36139 34901
rect 36998 34892 37004 34904
rect 37056 34892 37062 34944
rect 37274 34892 37280 34944
rect 37332 34932 37338 34944
rect 38013 34935 38071 34941
rect 38013 34932 38025 34935
rect 37332 34904 38025 34932
rect 37332 34892 37338 34904
rect 38013 34901 38025 34904
rect 38059 34901 38071 34935
rect 38013 34895 38071 34901
rect 38930 34892 38936 34944
rect 38988 34932 38994 34944
rect 40218 34932 40224 34944
rect 38988 34904 40224 34932
rect 38988 34892 38994 34904
rect 40218 34892 40224 34904
rect 40276 34932 40282 34944
rect 41233 34935 41291 34941
rect 41233 34932 41245 34935
rect 40276 34904 41245 34932
rect 40276 34892 40282 34904
rect 41233 34901 41245 34904
rect 41279 34901 41291 34935
rect 41233 34895 41291 34901
rect 45186 34892 45192 34944
rect 45244 34932 45250 34944
rect 46124 34941 46152 34972
rect 46998 34969 47010 34972
rect 47044 34969 47056 35003
rect 46998 34963 47056 34969
rect 45373 34935 45431 34941
rect 45373 34932 45385 34935
rect 45244 34904 45385 34932
rect 45244 34892 45250 34904
rect 45373 34901 45385 34904
rect 45419 34901 45431 34935
rect 45373 34895 45431 34901
rect 46109 34935 46167 34941
rect 46109 34901 46121 34935
rect 46155 34901 46167 34935
rect 46109 34895 46167 34901
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 25406 34688 25412 34740
rect 25464 34728 25470 34740
rect 25777 34731 25835 34737
rect 25777 34728 25789 34731
rect 25464 34700 25789 34728
rect 25464 34688 25470 34700
rect 25777 34697 25789 34700
rect 25823 34728 25835 34731
rect 25866 34728 25872 34740
rect 25823 34700 25872 34728
rect 25823 34697 25835 34700
rect 25777 34691 25835 34697
rect 25866 34688 25872 34700
rect 25924 34688 25930 34740
rect 26142 34688 26148 34740
rect 26200 34728 26206 34740
rect 27433 34731 27491 34737
rect 26200 34688 26234 34728
rect 27433 34697 27445 34731
rect 27479 34728 27491 34731
rect 27982 34728 27988 34740
rect 27479 34700 27988 34728
rect 27479 34697 27491 34700
rect 27433 34691 27491 34697
rect 27982 34688 27988 34700
rect 28040 34688 28046 34740
rect 32858 34728 32864 34740
rect 32819 34700 32864 34728
rect 32858 34688 32864 34700
rect 32916 34688 32922 34740
rect 33505 34731 33563 34737
rect 33505 34697 33517 34731
rect 33551 34728 33563 34731
rect 34882 34728 34888 34740
rect 33551 34700 34888 34728
rect 33551 34697 33563 34700
rect 33505 34691 33563 34697
rect 34882 34688 34888 34700
rect 34940 34688 34946 34740
rect 35894 34688 35900 34740
rect 35952 34728 35958 34740
rect 37553 34731 37611 34737
rect 37553 34728 37565 34731
rect 35952 34700 37565 34728
rect 35952 34688 35958 34700
rect 37553 34697 37565 34700
rect 37599 34697 37611 34731
rect 37553 34691 37611 34697
rect 39393 34731 39451 34737
rect 39393 34697 39405 34731
rect 39439 34728 39451 34731
rect 39942 34728 39948 34740
rect 39439 34700 39948 34728
rect 39439 34697 39451 34700
rect 39393 34691 39451 34697
rect 39942 34688 39948 34700
rect 40000 34688 40006 34740
rect 45373 34731 45431 34737
rect 45373 34697 45385 34731
rect 45419 34728 45431 34731
rect 45738 34728 45744 34740
rect 45419 34700 45744 34728
rect 45419 34697 45431 34700
rect 45373 34691 45431 34697
rect 45738 34688 45744 34700
rect 45796 34688 45802 34740
rect 46842 34728 46848 34740
rect 46803 34700 46848 34728
rect 46842 34688 46848 34700
rect 46900 34688 46906 34740
rect 26206 34660 26234 34688
rect 27249 34663 27307 34669
rect 27249 34660 27261 34663
rect 26206 34632 27261 34660
rect 27249 34629 27261 34632
rect 27295 34629 27307 34663
rect 27249 34623 27307 34629
rect 27522 34620 27528 34672
rect 27580 34660 27586 34672
rect 28138 34663 28196 34669
rect 28138 34660 28150 34663
rect 27580 34632 28150 34660
rect 27580 34620 27586 34632
rect 28138 34629 28150 34632
rect 28184 34629 28196 34663
rect 28138 34623 28196 34629
rect 29362 34620 29368 34672
rect 29420 34660 29426 34672
rect 29978 34663 30036 34669
rect 29978 34660 29990 34663
rect 29420 34632 29990 34660
rect 29420 34620 29426 34632
rect 29978 34629 29990 34632
rect 30024 34629 30036 34663
rect 34606 34660 34612 34672
rect 29978 34623 30036 34629
rect 34256 34632 34612 34660
rect 2038 34592 2044 34604
rect 1999 34564 2044 34592
rect 2038 34552 2044 34564
rect 2096 34552 2102 34604
rect 24394 34592 24400 34604
rect 24355 34564 24400 34592
rect 24394 34552 24400 34564
rect 24452 34552 24458 34604
rect 24486 34552 24492 34604
rect 24544 34592 24550 34604
rect 24653 34595 24711 34601
rect 24653 34592 24665 34595
rect 24544 34564 24665 34592
rect 24544 34552 24550 34564
rect 24653 34561 24665 34564
rect 24699 34561 24711 34595
rect 27062 34592 27068 34604
rect 27023 34564 27068 34592
rect 24653 34555 24711 34561
rect 27062 34552 27068 34564
rect 27120 34552 27126 34604
rect 27890 34592 27896 34604
rect 27851 34564 27896 34592
rect 27890 34552 27896 34564
rect 27948 34552 27954 34604
rect 32122 34592 32128 34604
rect 32083 34564 32128 34592
rect 32122 34552 32128 34564
rect 32180 34552 32186 34604
rect 32306 34592 32312 34604
rect 32267 34564 32312 34592
rect 32306 34552 32312 34564
rect 32364 34552 32370 34604
rect 32674 34592 32680 34604
rect 32635 34564 32680 34592
rect 32674 34552 32680 34564
rect 32732 34552 32738 34604
rect 33410 34592 33416 34604
rect 33371 34564 33416 34592
rect 33410 34552 33416 34564
rect 33468 34552 33474 34604
rect 33502 34552 33508 34604
rect 33560 34592 33566 34604
rect 34256 34601 34284 34632
rect 34606 34620 34612 34632
rect 34664 34620 34670 34672
rect 43806 34620 43812 34672
rect 43864 34660 43870 34672
rect 47762 34660 47768 34672
rect 43864 34632 47768 34660
rect 43864 34620 43870 34632
rect 33597 34595 33655 34601
rect 33597 34592 33609 34595
rect 33560 34564 33609 34592
rect 33560 34552 33566 34564
rect 33597 34561 33609 34564
rect 33643 34561 33655 34595
rect 33597 34555 33655 34561
rect 34241 34595 34299 34601
rect 34241 34561 34253 34595
rect 34287 34561 34299 34595
rect 34422 34592 34428 34604
rect 34383 34564 34428 34592
rect 34241 34555 34299 34561
rect 34422 34552 34428 34564
rect 34480 34552 34486 34604
rect 34514 34552 34520 34604
rect 34572 34592 34578 34604
rect 34572 34564 34617 34592
rect 34572 34552 34578 34564
rect 34698 34552 34704 34604
rect 34756 34592 34762 34604
rect 34974 34592 34980 34604
rect 34756 34564 34980 34592
rect 34756 34552 34762 34564
rect 34974 34552 34980 34564
rect 35032 34552 35038 34604
rect 35161 34595 35219 34601
rect 35161 34561 35173 34595
rect 35207 34592 35219 34595
rect 35342 34592 35348 34604
rect 35207 34564 35348 34592
rect 35207 34561 35219 34564
rect 35161 34555 35219 34561
rect 35342 34552 35348 34564
rect 35400 34552 35406 34604
rect 35621 34595 35679 34601
rect 35621 34561 35633 34595
rect 35667 34592 35679 34595
rect 35986 34592 35992 34604
rect 35667 34564 35992 34592
rect 35667 34561 35679 34564
rect 35621 34555 35679 34561
rect 35986 34552 35992 34564
rect 36044 34592 36050 34604
rect 36541 34595 36599 34601
rect 36541 34592 36553 34595
rect 36044 34564 36553 34592
rect 36044 34552 36050 34564
rect 36541 34561 36553 34564
rect 36587 34592 36599 34595
rect 36998 34592 37004 34604
rect 36587 34564 37004 34592
rect 36587 34561 36599 34564
rect 36541 34555 36599 34561
rect 36998 34552 37004 34564
rect 37056 34552 37062 34604
rect 37274 34592 37280 34604
rect 37235 34564 37280 34592
rect 37274 34552 37280 34564
rect 37332 34552 37338 34604
rect 37366 34552 37372 34604
rect 37424 34592 37430 34604
rect 39022 34592 39028 34604
rect 37424 34564 37469 34592
rect 38983 34564 39028 34592
rect 37424 34552 37430 34564
rect 39022 34552 39028 34564
rect 39080 34552 39086 34604
rect 41138 34592 41144 34604
rect 41099 34564 41144 34592
rect 41138 34552 41144 34564
rect 41196 34552 41202 34604
rect 42794 34552 42800 34604
rect 42852 34592 42858 34604
rect 43993 34595 44051 34601
rect 43993 34592 44005 34595
rect 42852 34564 44005 34592
rect 42852 34552 42858 34564
rect 43993 34561 44005 34564
rect 44039 34561 44051 34595
rect 43993 34555 44051 34561
rect 44260 34595 44318 34601
rect 44260 34561 44272 34595
rect 44306 34592 44318 34595
rect 45002 34592 45008 34604
rect 44306 34564 45008 34592
rect 44306 34561 44318 34564
rect 44260 34555 44318 34561
rect 45002 34552 45008 34564
rect 45060 34552 45066 34604
rect 46382 34552 46388 34604
rect 46440 34592 46446 34604
rect 46676 34601 46704 34632
rect 47762 34620 47768 34632
rect 47820 34620 47826 34672
rect 46477 34595 46535 34601
rect 46477 34592 46489 34595
rect 46440 34564 46489 34592
rect 46440 34552 46446 34564
rect 46477 34561 46489 34564
rect 46523 34561 46535 34595
rect 46477 34555 46535 34561
rect 46661 34595 46719 34601
rect 46661 34561 46673 34595
rect 46707 34561 46719 34595
rect 46661 34555 46719 34561
rect 2222 34524 2228 34536
rect 2183 34496 2228 34524
rect 2222 34484 2228 34496
rect 2280 34484 2286 34536
rect 3602 34524 3608 34536
rect 3563 34496 3608 34524
rect 3602 34484 3608 34496
rect 3660 34484 3666 34536
rect 29730 34524 29736 34536
rect 29691 34496 29736 34524
rect 29730 34484 29736 34496
rect 29788 34484 29794 34536
rect 32401 34527 32459 34533
rect 32401 34493 32413 34527
rect 32447 34493 32459 34527
rect 32401 34487 32459 34493
rect 32493 34527 32551 34533
rect 32493 34493 32505 34527
rect 32539 34493 32551 34527
rect 32493 34487 32551 34493
rect 32122 34416 32128 34468
rect 32180 34456 32186 34468
rect 32416 34456 32444 34487
rect 32180 34428 32444 34456
rect 32508 34456 32536 34487
rect 33962 34484 33968 34536
rect 34020 34524 34026 34536
rect 35713 34527 35771 34533
rect 35713 34524 35725 34527
rect 34020 34496 35725 34524
rect 34020 34484 34026 34496
rect 35713 34493 35725 34496
rect 35759 34493 35771 34527
rect 35713 34487 35771 34493
rect 36725 34527 36783 34533
rect 36725 34493 36737 34527
rect 36771 34524 36783 34527
rect 37384 34524 37412 34552
rect 36771 34496 37412 34524
rect 37553 34527 37611 34533
rect 36771 34493 36783 34496
rect 36725 34487 36783 34493
rect 37553 34493 37565 34527
rect 37599 34524 37611 34527
rect 38562 34524 38568 34536
rect 37599 34496 38568 34524
rect 37599 34493 37611 34496
rect 37553 34487 37611 34493
rect 32950 34456 32956 34468
rect 32508 34428 32956 34456
rect 32180 34416 32186 34428
rect 32950 34416 32956 34428
rect 33008 34456 33014 34468
rect 36740 34456 36768 34487
rect 38562 34484 38568 34496
rect 38620 34484 38626 34536
rect 39114 34524 39120 34536
rect 39075 34496 39120 34524
rect 39114 34484 39120 34496
rect 39172 34484 39178 34536
rect 41233 34527 41291 34533
rect 41233 34493 41245 34527
rect 41279 34524 41291 34527
rect 41690 34524 41696 34536
rect 41279 34496 41696 34524
rect 41279 34493 41291 34496
rect 41233 34487 41291 34493
rect 41690 34484 41696 34496
rect 41748 34484 41754 34536
rect 33008 34428 36768 34456
rect 33008 34416 33014 34428
rect 29270 34388 29276 34400
rect 29231 34360 29276 34388
rect 29270 34348 29276 34360
rect 29328 34348 29334 34400
rect 31110 34388 31116 34400
rect 31071 34360 31116 34388
rect 31110 34348 31116 34360
rect 31168 34348 31174 34400
rect 33318 34348 33324 34400
rect 33376 34388 33382 34400
rect 34057 34391 34115 34397
rect 34057 34388 34069 34391
rect 33376 34360 34069 34388
rect 33376 34348 33382 34360
rect 34057 34357 34069 34360
rect 34103 34357 34115 34391
rect 34057 34351 34115 34357
rect 34790 34348 34796 34400
rect 34848 34388 34854 34400
rect 35069 34391 35127 34397
rect 35069 34388 35081 34391
rect 34848 34360 35081 34388
rect 34848 34348 34854 34360
rect 35069 34357 35081 34360
rect 35115 34357 35127 34391
rect 35069 34351 35127 34357
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 2222 34144 2228 34196
rect 2280 34184 2286 34196
rect 2409 34187 2467 34193
rect 2409 34184 2421 34187
rect 2280 34156 2421 34184
rect 2280 34144 2286 34156
rect 2409 34153 2421 34156
rect 2455 34153 2467 34187
rect 2409 34147 2467 34153
rect 23661 34187 23719 34193
rect 23661 34153 23673 34187
rect 23707 34184 23719 34187
rect 24486 34184 24492 34196
rect 23707 34156 24492 34184
rect 23707 34153 23719 34156
rect 23661 34147 23719 34153
rect 24486 34144 24492 34156
rect 24544 34144 24550 34196
rect 27525 34187 27583 34193
rect 27525 34153 27537 34187
rect 27571 34184 27583 34187
rect 27614 34184 27620 34196
rect 27571 34156 27620 34184
rect 27571 34153 27583 34156
rect 27525 34147 27583 34153
rect 27614 34144 27620 34156
rect 27672 34184 27678 34196
rect 27890 34184 27896 34196
rect 27672 34156 27896 34184
rect 27672 34144 27678 34156
rect 27890 34144 27896 34156
rect 27948 34144 27954 34196
rect 31297 34187 31355 34193
rect 31297 34153 31309 34187
rect 31343 34184 31355 34187
rect 32306 34184 32312 34196
rect 31343 34156 32312 34184
rect 31343 34153 31355 34156
rect 31297 34147 31355 34153
rect 32306 34144 32312 34156
rect 32364 34144 32370 34196
rect 33229 34187 33287 34193
rect 33229 34184 33241 34187
rect 32508 34156 33241 34184
rect 32122 34116 32128 34128
rect 32083 34088 32128 34116
rect 32122 34076 32128 34088
rect 32180 34076 32186 34128
rect 32508 34057 32536 34156
rect 33229 34153 33241 34156
rect 33275 34153 33287 34187
rect 33229 34147 33287 34153
rect 36170 34144 36176 34196
rect 36228 34184 36234 34196
rect 36633 34187 36691 34193
rect 36633 34184 36645 34187
rect 36228 34156 36645 34184
rect 36228 34144 36234 34156
rect 36633 34153 36645 34156
rect 36679 34153 36691 34187
rect 36633 34147 36691 34153
rect 40862 34144 40868 34196
rect 40920 34184 40926 34196
rect 41049 34187 41107 34193
rect 41049 34184 41061 34187
rect 40920 34156 41061 34184
rect 40920 34144 40926 34156
rect 41049 34153 41061 34156
rect 41095 34153 41107 34187
rect 43806 34184 43812 34196
rect 43767 34156 43812 34184
rect 41049 34147 41107 34153
rect 43806 34144 43812 34156
rect 43864 34144 43870 34196
rect 45002 34184 45008 34196
rect 44963 34156 45008 34184
rect 45002 34144 45008 34156
rect 45060 34144 45066 34196
rect 33410 34116 33416 34128
rect 33152 34088 33416 34116
rect 24949 34051 25007 34057
rect 24949 34048 24961 34051
rect 23860 34020 24961 34048
rect 2317 33983 2375 33989
rect 2317 33949 2329 33983
rect 2363 33980 2375 33983
rect 2406 33980 2412 33992
rect 2363 33952 2412 33980
rect 2363 33949 2375 33952
rect 2317 33943 2375 33949
rect 2406 33940 2412 33952
rect 2464 33980 2470 33992
rect 18138 33980 18144 33992
rect 2464 33952 18144 33980
rect 2464 33940 2470 33952
rect 18138 33940 18144 33952
rect 18196 33940 18202 33992
rect 23860 33989 23888 34020
rect 24949 34017 24961 34020
rect 24995 34017 25007 34051
rect 24949 34011 25007 34017
rect 30745 34051 30803 34057
rect 30745 34017 30757 34051
rect 30791 34048 30803 34051
rect 32401 34051 32459 34057
rect 32401 34048 32413 34051
rect 30791 34020 31616 34048
rect 30791 34017 30803 34020
rect 30745 34011 30803 34017
rect 23845 33983 23903 33989
rect 23845 33949 23857 33983
rect 23891 33949 23903 33983
rect 23845 33943 23903 33949
rect 24673 33983 24731 33989
rect 24673 33949 24685 33983
rect 24719 33949 24731 33983
rect 24673 33943 24731 33949
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33980 24823 33983
rect 24854 33980 24860 33992
rect 24811 33952 24860 33980
rect 24811 33949 24823 33952
rect 24765 33943 24823 33949
rect 24688 33912 24716 33943
rect 24854 33940 24860 33952
rect 24912 33940 24918 33992
rect 29733 33983 29791 33989
rect 29733 33949 29745 33983
rect 29779 33980 29791 33983
rect 30374 33980 30380 33992
rect 29779 33952 30380 33980
rect 29779 33949 29791 33952
rect 29733 33943 29791 33949
rect 30374 33940 30380 33952
rect 30432 33940 30438 33992
rect 30650 33980 30656 33992
rect 30611 33952 30656 33980
rect 30650 33940 30656 33952
rect 30708 33940 30714 33992
rect 30837 33983 30895 33989
rect 30837 33949 30849 33983
rect 30883 33980 30895 33983
rect 31018 33980 31024 33992
rect 30883 33952 31024 33980
rect 30883 33949 30895 33952
rect 30837 33943 30895 33949
rect 31018 33940 31024 33952
rect 31076 33940 31082 33992
rect 31588 33989 31616 34020
rect 32140 34020 32413 34048
rect 32140 33992 32168 34020
rect 32401 34017 32413 34020
rect 32447 34017 32459 34051
rect 32401 34011 32459 34017
rect 32493 34051 32551 34057
rect 32493 34017 32505 34051
rect 32539 34017 32551 34051
rect 32493 34011 32551 34017
rect 31573 33983 31631 33989
rect 31573 33949 31585 33983
rect 31619 33980 31631 33983
rect 32122 33980 32128 33992
rect 31619 33952 32128 33980
rect 31619 33949 31631 33952
rect 31573 33943 31631 33949
rect 32122 33940 32128 33952
rect 32180 33940 32186 33992
rect 32214 33940 32220 33992
rect 32272 33980 32278 33992
rect 32309 33983 32367 33989
rect 32309 33980 32321 33983
rect 32272 33952 32321 33980
rect 32272 33940 32278 33952
rect 32309 33949 32321 33952
rect 32355 33949 32367 33983
rect 32309 33943 32367 33949
rect 25958 33912 25964 33924
rect 24688 33884 25964 33912
rect 25958 33872 25964 33884
rect 26016 33872 26022 33924
rect 26053 33915 26111 33921
rect 26053 33881 26065 33915
rect 26099 33912 26111 33915
rect 28626 33912 28632 33924
rect 26099 33884 28632 33912
rect 26099 33881 26111 33884
rect 26053 33875 26111 33881
rect 28626 33872 28632 33884
rect 28684 33872 28690 33924
rect 31297 33915 31355 33921
rect 31297 33881 31309 33915
rect 31343 33881 31355 33915
rect 31297 33875 31355 33881
rect 31481 33915 31539 33921
rect 31481 33881 31493 33915
rect 31527 33912 31539 33915
rect 32508 33912 32536 34011
rect 33152 33989 33180 34088
rect 33410 34076 33416 34088
rect 33468 34076 33474 34128
rect 36449 34051 36507 34057
rect 36449 34017 36461 34051
rect 36495 34048 36507 34051
rect 37918 34048 37924 34060
rect 36495 34020 37924 34048
rect 36495 34017 36507 34020
rect 36449 34011 36507 34017
rect 37918 34008 37924 34020
rect 37976 34008 37982 34060
rect 41690 34048 41696 34060
rect 41651 34020 41696 34048
rect 41690 34008 41696 34020
rect 41748 34008 41754 34060
rect 43349 34051 43407 34057
rect 43349 34017 43361 34051
rect 43395 34048 43407 34051
rect 46474 34048 46480 34060
rect 43395 34020 46480 34048
rect 43395 34017 43407 34020
rect 43349 34011 43407 34017
rect 46474 34008 46480 34020
rect 46532 34008 46538 34060
rect 46750 34048 46756 34060
rect 46711 34020 46756 34048
rect 46750 34008 46756 34020
rect 46808 34008 46814 34060
rect 32585 33983 32643 33989
rect 32585 33949 32597 33983
rect 32631 33949 32643 33983
rect 32585 33943 32643 33949
rect 33137 33983 33195 33989
rect 33137 33949 33149 33983
rect 33183 33949 33195 33983
rect 33137 33943 33195 33949
rect 33321 33983 33379 33989
rect 33321 33949 33333 33983
rect 33367 33980 33379 33983
rect 33410 33980 33416 33992
rect 33367 33952 33416 33980
rect 33367 33949 33379 33952
rect 33321 33943 33379 33949
rect 31527 33884 32536 33912
rect 32600 33912 32628 33943
rect 33410 33940 33416 33952
rect 33468 33940 33474 33992
rect 33962 33980 33968 33992
rect 33923 33952 33968 33980
rect 33962 33940 33968 33952
rect 34020 33940 34026 33992
rect 34698 33980 34704 33992
rect 34659 33952 34704 33980
rect 34698 33940 34704 33952
rect 34756 33940 34762 33992
rect 36354 33980 36360 33992
rect 36315 33952 36360 33980
rect 36354 33940 36360 33952
rect 36412 33940 36418 33992
rect 40586 33940 40592 33992
rect 40644 33980 40650 33992
rect 40681 33983 40739 33989
rect 40681 33980 40693 33983
rect 40644 33952 40693 33980
rect 40644 33940 40650 33952
rect 40681 33949 40693 33952
rect 40727 33949 40739 33983
rect 40681 33943 40739 33949
rect 40865 33983 40923 33989
rect 40865 33949 40877 33983
rect 40911 33949 40923 33983
rect 40865 33943 40923 33949
rect 33980 33912 34008 33940
rect 32600 33884 34008 33912
rect 34149 33915 34207 33921
rect 31527 33881 31539 33884
rect 31481 33875 31539 33881
rect 34149 33881 34161 33915
rect 34195 33912 34207 33915
rect 34422 33912 34428 33924
rect 34195 33884 34428 33912
rect 34195 33881 34207 33884
rect 34149 33875 34207 33881
rect 28994 33804 29000 33856
rect 29052 33844 29058 33856
rect 29549 33847 29607 33853
rect 29549 33844 29561 33847
rect 29052 33816 29561 33844
rect 29052 33804 29058 33816
rect 29549 33813 29561 33816
rect 29595 33813 29607 33847
rect 31312 33844 31340 33875
rect 34422 33872 34428 33884
rect 34480 33872 34486 33924
rect 34514 33872 34520 33924
rect 34572 33912 34578 33924
rect 34882 33912 34888 33924
rect 34572 33884 34888 33912
rect 34572 33872 34578 33884
rect 34882 33872 34888 33884
rect 34940 33912 34946 33924
rect 35342 33912 35348 33924
rect 34940 33884 35348 33912
rect 34940 33872 34946 33884
rect 35342 33872 35348 33884
rect 35400 33872 35406 33924
rect 40880 33912 40908 33943
rect 41230 33940 41236 33992
rect 41288 33980 41294 33992
rect 41509 33983 41567 33989
rect 41509 33980 41521 33983
rect 41288 33952 41521 33980
rect 41288 33940 41294 33952
rect 41509 33949 41521 33952
rect 41555 33949 41567 33983
rect 41509 33943 41567 33949
rect 42886 33940 42892 33992
rect 42944 33980 42950 33992
rect 43990 33980 43996 33992
rect 42944 33952 43996 33980
rect 42944 33940 42950 33952
rect 43990 33940 43996 33952
rect 44048 33940 44054 33992
rect 45186 33980 45192 33992
rect 45147 33952 45192 33980
rect 45186 33940 45192 33952
rect 45244 33940 45250 33992
rect 43254 33912 43260 33924
rect 40880 33884 43260 33912
rect 43254 33872 43260 33884
rect 43312 33872 43318 33924
rect 47020 33915 47078 33921
rect 47020 33881 47032 33915
rect 47066 33912 47078 33915
rect 47670 33912 47676 33924
rect 47066 33884 47676 33912
rect 47066 33881 47078 33884
rect 47020 33875 47078 33881
rect 47670 33872 47676 33884
rect 47728 33872 47734 33924
rect 32214 33844 32220 33856
rect 31312 33816 32220 33844
rect 29549 33807 29607 33813
rect 32214 33804 32220 33816
rect 32272 33804 32278 33856
rect 35066 33844 35072 33856
rect 35027 33816 35072 33844
rect 35066 33804 35072 33816
rect 35124 33804 35130 33856
rect 48038 33804 48044 33856
rect 48096 33844 48102 33856
rect 48133 33847 48191 33853
rect 48133 33844 48145 33847
rect 48096 33816 48145 33844
rect 48096 33804 48102 33816
rect 48133 33813 48145 33816
rect 48179 33813 48191 33847
rect 48133 33807 48191 33813
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 24394 33600 24400 33652
rect 24452 33600 24458 33652
rect 25498 33640 25504 33652
rect 25459 33612 25504 33640
rect 25498 33600 25504 33612
rect 25556 33600 25562 33652
rect 25961 33643 26019 33649
rect 25961 33609 25973 33643
rect 26007 33609 26019 33643
rect 25961 33603 26019 33609
rect 24412 33572 24440 33600
rect 24136 33544 24440 33572
rect 24136 33513 24164 33544
rect 24121 33507 24179 33513
rect 24121 33473 24133 33507
rect 24167 33473 24179 33507
rect 24121 33467 24179 33473
rect 24388 33507 24446 33513
rect 24388 33473 24400 33507
rect 24434 33504 24446 33507
rect 25976 33504 26004 33603
rect 31202 33600 31208 33652
rect 31260 33640 31266 33652
rect 34701 33643 34759 33649
rect 31260 33612 34652 33640
rect 31260 33600 31266 33612
rect 30926 33572 30932 33584
rect 30887 33544 30932 33572
rect 30926 33532 30932 33544
rect 30984 33532 30990 33584
rect 31018 33532 31024 33584
rect 31076 33572 31082 33584
rect 31076 33544 32536 33572
rect 31076 33532 31082 33544
rect 26142 33504 26148 33516
rect 24434 33476 26004 33504
rect 26103 33476 26148 33504
rect 24434 33473 24446 33476
rect 24388 33467 24446 33473
rect 26142 33464 26148 33476
rect 26200 33464 26206 33516
rect 28626 33504 28632 33516
rect 28539 33476 28632 33504
rect 28626 33464 28632 33476
rect 28684 33464 28690 33516
rect 31113 33507 31171 33513
rect 31113 33473 31125 33507
rect 31159 33504 31171 33507
rect 31202 33504 31208 33516
rect 31159 33476 31208 33504
rect 31159 33473 31171 33476
rect 31113 33467 31171 33473
rect 31202 33464 31208 33476
rect 31260 33464 31266 33516
rect 31662 33464 31668 33516
rect 31720 33504 31726 33516
rect 32508 33513 32536 33544
rect 33134 33532 33140 33584
rect 33192 33572 33198 33584
rect 33229 33575 33287 33581
rect 33229 33572 33241 33575
rect 33192 33544 33241 33572
rect 33192 33532 33198 33544
rect 33229 33541 33241 33544
rect 33275 33541 33287 33575
rect 34333 33575 34391 33581
rect 34333 33572 34345 33575
rect 33229 33535 33287 33541
rect 33704 33544 34345 33572
rect 33704 33516 33732 33544
rect 34333 33541 34345 33544
rect 34379 33541 34391 33575
rect 34624 33572 34652 33612
rect 34701 33609 34713 33643
rect 34747 33640 34759 33643
rect 35066 33640 35072 33652
rect 34747 33612 35072 33640
rect 34747 33609 34759 33612
rect 34701 33603 34759 33609
rect 35066 33600 35072 33612
rect 35124 33600 35130 33652
rect 41230 33640 41236 33652
rect 41191 33612 41236 33640
rect 41230 33600 41236 33612
rect 41288 33600 41294 33652
rect 43254 33600 43260 33652
rect 43312 33640 43318 33652
rect 46845 33643 46903 33649
rect 46845 33640 46857 33643
rect 43312 33612 46857 33640
rect 43312 33600 43318 33612
rect 46845 33609 46857 33612
rect 46891 33609 46903 33643
rect 46845 33603 46903 33609
rect 42886 33572 42892 33584
rect 34624 33544 42892 33572
rect 34333 33535 34391 33541
rect 42886 33532 42892 33544
rect 42944 33532 42950 33584
rect 43064 33575 43122 33581
rect 43064 33541 43076 33575
rect 43110 33572 43122 33575
rect 43438 33572 43444 33584
rect 43110 33544 43444 33572
rect 43110 33541 43122 33544
rect 43064 33535 43122 33541
rect 43438 33532 43444 33544
rect 43496 33532 43502 33584
rect 32401 33507 32459 33513
rect 32401 33504 32413 33507
rect 31720 33476 32413 33504
rect 31720 33464 31726 33476
rect 32401 33473 32413 33476
rect 32447 33473 32459 33507
rect 32401 33467 32459 33473
rect 32493 33507 32551 33513
rect 32493 33473 32505 33507
rect 32539 33504 32551 33507
rect 33318 33504 33324 33516
rect 32539 33476 33324 33504
rect 32539 33473 32551 33476
rect 32493 33467 32551 33473
rect 33318 33464 33324 33476
rect 33376 33464 33382 33516
rect 33502 33504 33508 33516
rect 33463 33476 33508 33504
rect 33502 33464 33508 33476
rect 33560 33464 33566 33516
rect 33594 33507 33652 33513
rect 33594 33473 33606 33507
rect 33640 33473 33652 33507
rect 33594 33467 33652 33473
rect 33689 33510 33747 33516
rect 33689 33476 33701 33510
rect 33735 33476 33747 33510
rect 33689 33470 33747 33476
rect 28644 33368 28672 33464
rect 29730 33396 29736 33448
rect 29788 33436 29794 33448
rect 30285 33439 30343 33445
rect 30285 33436 30297 33439
rect 29788 33408 30297 33436
rect 29788 33396 29794 33408
rect 30285 33405 30297 33408
rect 30331 33436 30343 33439
rect 31754 33436 31760 33448
rect 30331 33408 31760 33436
rect 30331 33405 30343 33408
rect 30285 33399 30343 33405
rect 31754 33396 31760 33408
rect 31812 33396 31818 33448
rect 32214 33396 32220 33448
rect 32272 33436 32278 33448
rect 32309 33439 32367 33445
rect 32309 33436 32321 33439
rect 32272 33408 32321 33436
rect 32272 33396 32278 33408
rect 32309 33405 32321 33408
rect 32355 33405 32367 33439
rect 32309 33399 32367 33405
rect 32582 33396 32588 33448
rect 32640 33436 32646 33448
rect 32640 33408 32685 33436
rect 32640 33396 32646 33408
rect 33042 33396 33048 33448
rect 33100 33436 33106 33448
rect 33609 33436 33637 33467
rect 33870 33464 33876 33516
rect 33928 33504 33934 33516
rect 33928 33476 33973 33504
rect 33928 33464 33934 33476
rect 34422 33464 34428 33516
rect 34480 33504 34486 33516
rect 34517 33507 34575 33513
rect 34517 33504 34529 33507
rect 34480 33476 34529 33504
rect 34480 33464 34486 33476
rect 34517 33473 34529 33476
rect 34563 33473 34575 33507
rect 34790 33504 34796 33516
rect 34751 33476 34796 33504
rect 34517 33467 34575 33473
rect 34790 33464 34796 33476
rect 34848 33464 34854 33516
rect 41414 33464 41420 33516
rect 41472 33504 41478 33516
rect 42794 33504 42800 33516
rect 41472 33476 41517 33504
rect 42755 33476 42800 33504
rect 41472 33464 41478 33476
rect 42794 33464 42800 33476
rect 42852 33464 42858 33516
rect 44818 33504 44824 33516
rect 44779 33476 44824 33504
rect 44818 33464 44824 33476
rect 44876 33464 44882 33516
rect 46842 33464 46848 33516
rect 46900 33504 46906 33516
rect 47029 33507 47087 33513
rect 47029 33504 47041 33507
rect 46900 33476 47041 33504
rect 46900 33464 46906 33476
rect 47029 33473 47041 33476
rect 47075 33473 47087 33507
rect 47029 33467 47087 33473
rect 33100 33408 33637 33436
rect 33100 33396 33106 33408
rect 38102 33368 38108 33380
rect 28644 33340 38108 33368
rect 38102 33328 38108 33340
rect 38160 33328 38166 33380
rect 44177 33371 44235 33377
rect 44177 33337 44189 33371
rect 44223 33368 44235 33371
rect 44726 33368 44732 33380
rect 44223 33340 44732 33368
rect 44223 33337 44235 33340
rect 44177 33331 44235 33337
rect 44726 33328 44732 33340
rect 44784 33328 44790 33380
rect 32125 33303 32183 33309
rect 32125 33269 32137 33303
rect 32171 33300 32183 33303
rect 32490 33300 32496 33312
rect 32171 33272 32496 33300
rect 32171 33269 32183 33272
rect 32125 33263 32183 33269
rect 32490 33260 32496 33272
rect 32548 33260 32554 33312
rect 33226 33260 33232 33312
rect 33284 33300 33290 33312
rect 35802 33300 35808 33312
rect 33284 33272 35808 33300
rect 33284 33260 33290 33272
rect 35802 33260 35808 33272
rect 35860 33260 35866 33312
rect 44634 33300 44640 33312
rect 44595 33272 44640 33300
rect 44634 33260 44640 33272
rect 44692 33260 44698 33312
rect 46934 33260 46940 33312
rect 46992 33300 46998 33312
rect 47765 33303 47823 33309
rect 47765 33300 47777 33303
rect 46992 33272 47777 33300
rect 46992 33260 46998 33272
rect 47765 33269 47777 33272
rect 47811 33269 47823 33303
rect 47765 33263 47823 33269
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 24857 33099 24915 33105
rect 24857 33065 24869 33099
rect 24903 33096 24915 33099
rect 26142 33096 26148 33108
rect 24903 33068 26148 33096
rect 24903 33065 24915 33068
rect 24857 33059 24915 33065
rect 26142 33056 26148 33068
rect 26200 33056 26206 33108
rect 30374 33096 30380 33108
rect 30335 33068 30380 33096
rect 30374 33056 30380 33068
rect 30432 33056 30438 33108
rect 30650 33056 30656 33108
rect 30708 33096 30714 33108
rect 31662 33096 31668 33108
rect 30708 33068 31668 33096
rect 30708 33056 30714 33068
rect 31662 33056 31668 33068
rect 31720 33056 31726 33108
rect 32582 33056 32588 33108
rect 32640 33096 32646 33108
rect 33045 33099 33103 33105
rect 33045 33096 33057 33099
rect 32640 33068 33057 33096
rect 32640 33056 32646 33068
rect 33045 33065 33057 33068
rect 33091 33065 33103 33099
rect 33045 33059 33103 33065
rect 33134 33056 33140 33108
rect 33192 33096 33198 33108
rect 33192 33068 36308 33096
rect 33192 33056 33198 33068
rect 32306 33028 32312 33040
rect 30208 33000 32312 33028
rect 24854 32960 24860 32972
rect 24688 32932 24860 32960
rect 2130 32852 2136 32904
rect 2188 32892 2194 32904
rect 24688 32901 24716 32932
rect 24854 32920 24860 32932
rect 24912 32960 24918 32972
rect 27614 32960 27620 32972
rect 24912 32932 25544 32960
rect 27575 32932 27620 32960
rect 24912 32920 24918 32932
rect 2317 32895 2375 32901
rect 2317 32892 2329 32895
rect 2188 32864 2329 32892
rect 2188 32852 2194 32864
rect 2317 32861 2329 32864
rect 2363 32861 2375 32895
rect 2317 32855 2375 32861
rect 24581 32895 24639 32901
rect 24581 32861 24593 32895
rect 24627 32861 24639 32895
rect 24581 32855 24639 32861
rect 24673 32895 24731 32901
rect 24673 32861 24685 32895
rect 24719 32861 24731 32895
rect 25406 32892 25412 32904
rect 25367 32864 25412 32892
rect 24673 32855 24731 32861
rect 24596 32824 24624 32855
rect 25406 32852 25412 32864
rect 25464 32852 25470 32904
rect 25516 32901 25544 32932
rect 27614 32920 27620 32932
rect 27672 32920 27678 32972
rect 29270 32920 29276 32972
rect 29328 32960 29334 32972
rect 29546 32960 29552 32972
rect 29328 32932 29552 32960
rect 29328 32920 29334 32932
rect 29546 32920 29552 32932
rect 29604 32960 29610 32972
rect 30009 32963 30067 32969
rect 30009 32960 30021 32963
rect 29604 32932 30021 32960
rect 29604 32920 29610 32932
rect 30009 32929 30021 32932
rect 30055 32929 30067 32963
rect 30009 32923 30067 32929
rect 25501 32895 25559 32901
rect 25501 32861 25513 32895
rect 25547 32892 25559 32895
rect 26329 32895 26387 32901
rect 25547 32864 26188 32892
rect 25547 32861 25559 32864
rect 25501 32855 25559 32861
rect 26050 32824 26056 32836
rect 24596 32796 26056 32824
rect 26050 32784 26056 32796
rect 26108 32784 26114 32836
rect 25314 32716 25320 32768
rect 25372 32756 25378 32768
rect 26160 32765 26188 32864
rect 26329 32861 26341 32895
rect 26375 32861 26387 32895
rect 26329 32855 26387 32861
rect 27884 32895 27942 32901
rect 27884 32861 27896 32895
rect 27930 32892 27942 32895
rect 28994 32892 29000 32904
rect 27930 32864 29000 32892
rect 27930 32861 27942 32864
rect 27884 32855 27942 32861
rect 26344 32824 26372 32855
rect 28994 32852 29000 32864
rect 29052 32852 29058 32904
rect 30208 32901 30236 33000
rect 32306 32988 32312 33000
rect 32364 32988 32370 33040
rect 32490 32988 32496 33040
rect 32548 33028 32554 33040
rect 34330 33028 34336 33040
rect 32548 33000 34336 33028
rect 32548 32988 32554 33000
rect 34330 32988 34336 33000
rect 34388 32988 34394 33040
rect 36280 33028 36308 33068
rect 36354 33056 36360 33108
rect 36412 33096 36418 33108
rect 37369 33099 37427 33105
rect 37369 33096 37381 33099
rect 36412 33068 37381 33096
rect 36412 33056 36418 33068
rect 37369 33065 37381 33068
rect 37415 33065 37427 33099
rect 37369 33059 37427 33065
rect 38654 33056 38660 33108
rect 38712 33096 38718 33108
rect 39758 33096 39764 33108
rect 38712 33068 39764 33096
rect 38712 33056 38718 33068
rect 39758 33056 39764 33068
rect 39816 33096 39822 33108
rect 40037 33099 40095 33105
rect 40037 33096 40049 33099
rect 39816 33068 40049 33096
rect 39816 33056 39822 33068
rect 40037 33065 40049 33068
rect 40083 33065 40095 33099
rect 40770 33096 40776 33108
rect 40731 33068 40776 33096
rect 40037 33059 40095 33065
rect 40770 33056 40776 33068
rect 40828 33056 40834 33108
rect 40957 33099 41015 33105
rect 40957 33065 40969 33099
rect 41003 33096 41015 33099
rect 41414 33096 41420 33108
rect 41003 33068 41420 33096
rect 41003 33065 41015 33068
rect 40957 33059 41015 33065
rect 41414 33056 41420 33068
rect 41472 33056 41478 33108
rect 42794 33056 42800 33108
rect 42852 33096 42858 33108
rect 42889 33099 42947 33105
rect 42889 33096 42901 33099
rect 42852 33068 42901 33096
rect 42852 33056 42858 33068
rect 42889 33065 42901 33068
rect 42935 33065 42947 33099
rect 42889 33059 42947 33065
rect 43809 33099 43867 33105
rect 43809 33065 43821 33099
rect 43855 33096 43867 33099
rect 44174 33096 44180 33108
rect 43855 33068 44180 33096
rect 43855 33065 43867 33068
rect 43809 33059 43867 33065
rect 40126 33028 40132 33040
rect 36280 33000 40132 33028
rect 40126 32988 40132 33000
rect 40184 33028 40190 33040
rect 41690 33028 41696 33040
rect 40184 33000 41696 33028
rect 40184 32988 40190 33000
rect 41690 32988 41696 33000
rect 41748 32988 41754 33040
rect 31389 32963 31447 32969
rect 31389 32929 31401 32963
rect 31435 32960 31447 32963
rect 35713 32963 35771 32969
rect 31435 32932 33272 32960
rect 31435 32929 31447 32932
rect 31389 32923 31447 32929
rect 33244 32904 33272 32932
rect 35713 32929 35725 32963
rect 35759 32960 35771 32963
rect 35894 32960 35900 32972
rect 35759 32932 35900 32960
rect 35759 32929 35771 32932
rect 35713 32923 35771 32929
rect 35894 32920 35900 32932
rect 35952 32960 35958 32972
rect 37093 32963 37151 32969
rect 37093 32960 37105 32963
rect 35952 32932 37105 32960
rect 35952 32920 35958 32932
rect 37093 32929 37105 32932
rect 37139 32960 37151 32963
rect 42904 32960 42932 33059
rect 44174 33056 44180 33068
rect 44232 33096 44238 33108
rect 47670 33096 47676 33108
rect 44232 33068 47072 33096
rect 47631 33068 47676 33096
rect 44232 33056 44238 33068
rect 45005 32963 45063 32969
rect 45005 32960 45017 32963
rect 37139 32932 38608 32960
rect 42904 32932 45017 32960
rect 37139 32929 37151 32932
rect 37093 32923 37151 32929
rect 30193 32895 30251 32901
rect 30193 32861 30205 32895
rect 30239 32861 30251 32895
rect 31294 32892 31300 32904
rect 31255 32864 31300 32892
rect 30193 32855 30251 32861
rect 31294 32852 31300 32864
rect 31352 32852 31358 32904
rect 32309 32895 32367 32901
rect 32309 32861 32321 32895
rect 32355 32861 32367 32895
rect 32309 32855 32367 32861
rect 30374 32824 30380 32836
rect 26344 32796 30380 32824
rect 30374 32784 30380 32796
rect 30432 32824 30438 32836
rect 31202 32824 31208 32836
rect 30432 32796 31208 32824
rect 30432 32784 30438 32796
rect 31202 32784 31208 32796
rect 31260 32784 31266 32836
rect 32324 32824 32352 32855
rect 32398 32852 32404 32904
rect 32456 32892 32462 32904
rect 32585 32895 32643 32901
rect 32585 32892 32597 32895
rect 32456 32864 32597 32892
rect 32456 32852 32462 32864
rect 32585 32861 32597 32864
rect 32631 32861 32643 32895
rect 33226 32892 33232 32904
rect 33187 32864 33232 32892
rect 32585 32855 32643 32861
rect 33226 32852 33232 32864
rect 33284 32852 33290 32904
rect 33410 32892 33416 32904
rect 33371 32864 33416 32892
rect 33410 32852 33416 32864
rect 33468 32852 33474 32904
rect 33505 32895 33563 32901
rect 33505 32861 33517 32895
rect 33551 32894 33563 32895
rect 35529 32895 35587 32901
rect 33551 32892 33732 32894
rect 33551 32866 33916 32892
rect 33551 32861 33563 32866
rect 33505 32855 33563 32861
rect 33134 32824 33140 32836
rect 32324 32796 33140 32824
rect 33134 32784 33140 32796
rect 33192 32784 33198 32836
rect 25685 32759 25743 32765
rect 25685 32756 25697 32759
rect 25372 32728 25697 32756
rect 25372 32716 25378 32728
rect 25685 32725 25697 32728
rect 25731 32725 25743 32759
rect 25685 32719 25743 32725
rect 26145 32759 26203 32765
rect 26145 32725 26157 32759
rect 26191 32725 26203 32759
rect 26145 32719 26203 32725
rect 28810 32716 28816 32768
rect 28868 32756 28874 32768
rect 28997 32759 29055 32765
rect 28997 32756 29009 32759
rect 28868 32728 29009 32756
rect 28868 32716 28874 32728
rect 28997 32725 29009 32728
rect 29043 32725 29055 32759
rect 28997 32719 29055 32725
rect 32125 32759 32183 32765
rect 32125 32725 32137 32759
rect 32171 32756 32183 32759
rect 32306 32756 32312 32768
rect 32171 32728 32312 32756
rect 32171 32725 32183 32728
rect 32125 32719 32183 32725
rect 32306 32716 32312 32728
rect 32364 32716 32370 32768
rect 32490 32756 32496 32768
rect 32451 32728 32496 32756
rect 32490 32716 32496 32728
rect 32548 32716 32554 32768
rect 32674 32716 32680 32768
rect 32732 32756 32738 32768
rect 33612 32756 33640 32866
rect 33704 32864 33916 32866
rect 33888 32824 33916 32864
rect 35529 32861 35541 32895
rect 35575 32892 35587 32895
rect 35802 32892 35808 32904
rect 35575 32864 35808 32892
rect 35575 32861 35587 32864
rect 35529 32855 35587 32861
rect 35802 32852 35808 32864
rect 35860 32852 35866 32904
rect 37001 32895 37059 32901
rect 37001 32861 37013 32895
rect 37047 32892 37059 32895
rect 37274 32892 37280 32904
rect 37047 32864 37280 32892
rect 37047 32861 37059 32864
rect 37001 32855 37059 32861
rect 37274 32852 37280 32864
rect 37332 32892 37338 32904
rect 38010 32892 38016 32904
rect 37332 32864 38016 32892
rect 37332 32852 37338 32864
rect 38010 32852 38016 32864
rect 38068 32852 38074 32904
rect 38580 32836 38608 32932
rect 45005 32929 45017 32932
rect 45051 32929 45063 32963
rect 45005 32923 45063 32929
rect 43990 32892 43996 32904
rect 43951 32864 43996 32892
rect 43990 32852 43996 32864
rect 44048 32852 44054 32904
rect 44634 32852 44640 32904
rect 44692 32892 44698 32904
rect 47044 32901 47072 33068
rect 47670 33056 47676 33068
rect 47728 33056 47734 33108
rect 45261 32895 45319 32901
rect 45261 32892 45273 32895
rect 44692 32864 45273 32892
rect 44692 32852 44698 32864
rect 45261 32861 45273 32864
rect 45307 32861 45319 32895
rect 46845 32895 46903 32901
rect 46845 32892 46857 32895
rect 45261 32855 45319 32861
rect 46400 32864 46857 32892
rect 35986 32824 35992 32836
rect 33888 32796 35992 32824
rect 35986 32784 35992 32796
rect 36044 32784 36050 32836
rect 38562 32784 38568 32836
rect 38620 32824 38626 32836
rect 39945 32827 40003 32833
rect 39945 32824 39957 32827
rect 38620 32796 39957 32824
rect 38620 32784 38626 32796
rect 39945 32793 39957 32796
rect 39991 32793 40003 32827
rect 39945 32787 40003 32793
rect 40589 32827 40647 32833
rect 40589 32793 40601 32827
rect 40635 32824 40647 32827
rect 40954 32824 40960 32836
rect 40635 32796 40960 32824
rect 40635 32793 40647 32796
rect 40589 32787 40647 32793
rect 40954 32784 40960 32796
rect 41012 32784 41018 32836
rect 41598 32824 41604 32836
rect 41559 32796 41604 32824
rect 41598 32784 41604 32796
rect 41656 32784 41662 32836
rect 32732 32728 33640 32756
rect 32732 32716 32738 32728
rect 40494 32716 40500 32768
rect 40552 32756 40558 32768
rect 40789 32759 40847 32765
rect 40789 32756 40801 32759
rect 40552 32728 40801 32756
rect 40552 32716 40558 32728
rect 40789 32725 40801 32728
rect 40835 32725 40847 32759
rect 40789 32719 40847 32725
rect 46106 32716 46112 32768
rect 46164 32756 46170 32768
rect 46400 32765 46428 32864
rect 46845 32861 46857 32864
rect 46891 32861 46903 32895
rect 46845 32855 46903 32861
rect 47029 32895 47087 32901
rect 47029 32861 47041 32895
rect 47075 32861 47087 32895
rect 47029 32855 47087 32861
rect 47213 32895 47271 32901
rect 47213 32861 47225 32895
rect 47259 32892 47271 32895
rect 47857 32895 47915 32901
rect 47857 32892 47869 32895
rect 47259 32864 47869 32892
rect 47259 32861 47271 32864
rect 47213 32855 47271 32861
rect 47857 32861 47869 32864
rect 47903 32861 47915 32895
rect 47857 32855 47915 32861
rect 47044 32824 47072 32855
rect 47302 32824 47308 32836
rect 47044 32796 47308 32824
rect 47302 32784 47308 32796
rect 47360 32784 47366 32836
rect 46385 32759 46443 32765
rect 46385 32756 46397 32759
rect 46164 32728 46397 32756
rect 46164 32716 46170 32728
rect 46385 32725 46397 32728
rect 46431 32725 46443 32759
rect 46385 32719 46443 32725
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 29546 32552 29552 32564
rect 28736 32524 29552 32552
rect 2130 32416 2136 32428
rect 2091 32388 2136 32416
rect 2130 32376 2136 32388
rect 2188 32376 2194 32428
rect 25314 32416 25320 32428
rect 25275 32388 25320 32416
rect 25314 32376 25320 32388
rect 25372 32376 25378 32428
rect 28537 32419 28595 32425
rect 28537 32385 28549 32419
rect 28583 32416 28595 32419
rect 28736 32416 28764 32524
rect 29546 32512 29552 32524
rect 29604 32512 29610 32564
rect 29730 32552 29736 32564
rect 29691 32524 29736 32552
rect 29730 32512 29736 32524
rect 29788 32512 29794 32564
rect 32490 32552 32496 32564
rect 32451 32524 32496 32552
rect 32490 32512 32496 32524
rect 32548 32512 32554 32564
rect 33134 32512 33140 32564
rect 33192 32552 33198 32564
rect 34422 32552 34428 32564
rect 33192 32524 34428 32552
rect 33192 32512 33198 32524
rect 34422 32512 34428 32524
rect 34480 32512 34486 32564
rect 35713 32555 35771 32561
rect 35713 32521 35725 32555
rect 35759 32552 35771 32555
rect 37090 32552 37096 32564
rect 35759 32524 37096 32552
rect 35759 32521 35771 32524
rect 35713 32515 35771 32521
rect 37090 32512 37096 32524
rect 37148 32552 37154 32564
rect 37277 32555 37335 32561
rect 37277 32552 37289 32555
rect 37148 32524 37289 32552
rect 37148 32512 37154 32524
rect 37277 32521 37289 32524
rect 37323 32521 37335 32555
rect 37918 32552 37924 32564
rect 37879 32524 37924 32552
rect 37277 32515 37335 32521
rect 37918 32512 37924 32524
rect 37976 32512 37982 32564
rect 38654 32552 38660 32564
rect 38028 32524 38660 32552
rect 28810 32444 28816 32496
rect 28868 32484 28874 32496
rect 28868 32456 29868 32484
rect 28868 32444 28874 32456
rect 28583 32388 28764 32416
rect 29022 32419 29080 32425
rect 28583 32385 28595 32388
rect 28537 32379 28595 32385
rect 29022 32385 29034 32419
rect 29068 32416 29080 32419
rect 29178 32416 29184 32428
rect 29068 32388 29184 32416
rect 29068 32385 29080 32388
rect 29022 32379 29080 32385
rect 29178 32376 29184 32388
rect 29236 32376 29242 32428
rect 29840 32425 29868 32456
rect 31662 32444 31668 32496
rect 31720 32484 31726 32496
rect 32125 32487 32183 32493
rect 32125 32484 32137 32487
rect 31720 32456 32137 32484
rect 31720 32444 31726 32456
rect 32125 32453 32137 32456
rect 32171 32453 32183 32487
rect 32125 32447 32183 32453
rect 32309 32487 32367 32493
rect 32309 32453 32321 32487
rect 32355 32484 32367 32487
rect 33318 32484 33324 32496
rect 32355 32456 33324 32484
rect 32355 32453 32367 32456
rect 32309 32447 32367 32453
rect 33318 32444 33324 32456
rect 33376 32444 33382 32496
rect 33410 32444 33416 32496
rect 33468 32484 33474 32496
rect 34146 32484 34152 32496
rect 33468 32456 34152 32484
rect 33468 32444 33474 32456
rect 34146 32444 34152 32456
rect 34204 32444 34210 32496
rect 34330 32444 34336 32496
rect 34388 32484 34394 32496
rect 36446 32484 36452 32496
rect 34388 32456 36452 32484
rect 34388 32444 34394 32456
rect 29641 32419 29699 32425
rect 29641 32385 29653 32419
rect 29687 32385 29699 32419
rect 29641 32379 29699 32385
rect 29825 32419 29883 32425
rect 29825 32385 29837 32419
rect 29871 32385 29883 32419
rect 30834 32416 30840 32428
rect 30795 32388 30840 32416
rect 29825 32379 29883 32385
rect 2317 32351 2375 32357
rect 2317 32317 2329 32351
rect 2363 32348 2375 32351
rect 2498 32348 2504 32360
rect 2363 32320 2504 32348
rect 2363 32317 2375 32320
rect 2317 32311 2375 32317
rect 2498 32308 2504 32320
rect 2556 32308 2562 32360
rect 2774 32348 2780 32360
rect 2735 32320 2780 32348
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 27614 32308 27620 32360
rect 27672 32348 27678 32360
rect 28810 32348 28816 32360
rect 27672 32320 28816 32348
rect 27672 32308 27678 32320
rect 28810 32308 28816 32320
rect 28868 32308 28874 32360
rect 28905 32351 28963 32357
rect 28905 32317 28917 32351
rect 28951 32348 28963 32351
rect 29656 32348 29684 32379
rect 30834 32376 30840 32388
rect 30892 32376 30898 32428
rect 35728 32425 35756 32456
rect 36446 32444 36452 32456
rect 36504 32484 36510 32496
rect 36504 32456 36584 32484
rect 36504 32444 36510 32456
rect 35529 32419 35587 32425
rect 35529 32385 35541 32419
rect 35575 32385 35587 32419
rect 35529 32379 35587 32385
rect 35713 32419 35771 32425
rect 35713 32385 35725 32419
rect 35759 32385 35771 32419
rect 36354 32416 36360 32428
rect 36315 32388 36360 32416
rect 35713 32379 35771 32385
rect 31110 32348 31116 32360
rect 28951 32320 31116 32348
rect 28951 32317 28963 32320
rect 28905 32311 28963 32317
rect 27798 32240 27804 32292
rect 27856 32280 27862 32292
rect 28920 32280 28948 32311
rect 31110 32308 31116 32320
rect 31168 32308 31174 32360
rect 35544 32348 35572 32379
rect 36354 32376 36360 32388
rect 36412 32376 36418 32428
rect 36556 32425 36584 32456
rect 36541 32419 36599 32425
rect 36541 32385 36553 32419
rect 36587 32385 36599 32419
rect 36541 32379 36599 32385
rect 37737 32419 37795 32425
rect 37737 32385 37749 32419
rect 37783 32416 37795 32419
rect 38028 32416 38056 32524
rect 38654 32512 38660 32524
rect 38712 32512 38718 32564
rect 39022 32512 39028 32564
rect 39080 32552 39086 32564
rect 39209 32555 39267 32561
rect 39209 32552 39221 32555
rect 39080 32524 39221 32552
rect 39080 32512 39086 32524
rect 39209 32521 39221 32524
rect 39255 32521 39267 32555
rect 39209 32515 39267 32521
rect 39577 32555 39635 32561
rect 39577 32521 39589 32555
rect 39623 32552 39635 32555
rect 40034 32552 40040 32564
rect 39623 32524 40040 32552
rect 39623 32521 39635 32524
rect 39577 32515 39635 32521
rect 40034 32512 40040 32524
rect 40092 32552 40098 32564
rect 40865 32555 40923 32561
rect 40865 32552 40877 32555
rect 40092 32524 40877 32552
rect 40092 32512 40098 32524
rect 40865 32521 40877 32524
rect 40911 32521 40923 32555
rect 40865 32515 40923 32521
rect 40954 32512 40960 32564
rect 41012 32552 41018 32564
rect 41417 32555 41475 32561
rect 41417 32552 41429 32555
rect 41012 32524 41429 32552
rect 41012 32512 41018 32524
rect 41417 32521 41429 32524
rect 41463 32521 41475 32555
rect 41417 32515 41475 32521
rect 43717 32555 43775 32561
rect 43717 32521 43729 32555
rect 43763 32552 43775 32555
rect 44818 32552 44824 32564
rect 43763 32524 44824 32552
rect 43763 32521 43775 32524
rect 43717 32515 43775 32521
rect 44818 32512 44824 32524
rect 44876 32512 44882 32564
rect 38672 32456 39712 32484
rect 38562 32416 38568 32428
rect 37783 32388 38056 32416
rect 38523 32388 38568 32416
rect 37783 32385 37795 32388
rect 37737 32379 37795 32385
rect 38562 32376 38568 32388
rect 38620 32376 38626 32428
rect 36170 32348 36176 32360
rect 35544 32320 36176 32348
rect 36170 32308 36176 32320
rect 36228 32348 36234 32360
rect 36449 32351 36507 32357
rect 36449 32348 36461 32351
rect 36228 32320 36461 32348
rect 36228 32308 36234 32320
rect 36449 32317 36461 32320
rect 36495 32317 36507 32351
rect 36449 32311 36507 32317
rect 36630 32308 36636 32360
rect 36688 32348 36694 32360
rect 37642 32348 37648 32360
rect 36688 32320 36733 32348
rect 37603 32320 37648 32348
rect 36688 32308 36694 32320
rect 37642 32308 37648 32320
rect 37700 32308 37706 32360
rect 38378 32348 38384 32360
rect 38339 32320 38384 32348
rect 38378 32308 38384 32320
rect 38436 32308 38442 32360
rect 29178 32280 29184 32292
rect 27856 32252 28948 32280
rect 29091 32252 29184 32280
rect 27856 32240 27862 32252
rect 29178 32240 29184 32252
rect 29236 32280 29242 32292
rect 30282 32280 30288 32292
rect 29236 32252 30288 32280
rect 29236 32240 29242 32252
rect 30282 32240 30288 32252
rect 30340 32240 30346 32292
rect 38672 32280 38700 32456
rect 39684 32425 39712 32456
rect 39758 32444 39764 32496
rect 39816 32484 39822 32496
rect 40221 32487 40279 32493
rect 39816 32456 40172 32484
rect 39816 32444 39822 32456
rect 39393 32419 39451 32425
rect 39393 32385 39405 32419
rect 39439 32385 39451 32419
rect 39393 32379 39451 32385
rect 39669 32419 39727 32425
rect 39669 32385 39681 32419
rect 39715 32416 39727 32419
rect 39942 32416 39948 32428
rect 39715 32388 39948 32416
rect 39715 32385 39727 32388
rect 39669 32379 39727 32385
rect 38749 32351 38807 32357
rect 38749 32317 38761 32351
rect 38795 32348 38807 32351
rect 39408 32348 39436 32379
rect 39942 32376 39948 32388
rect 40000 32376 40006 32428
rect 40144 32425 40172 32456
rect 40221 32453 40233 32487
rect 40267 32484 40279 32487
rect 40267 32456 41000 32484
rect 40267 32453 40279 32456
rect 40221 32447 40279 32453
rect 40129 32419 40187 32425
rect 40129 32385 40141 32419
rect 40175 32385 40187 32419
rect 40310 32416 40316 32428
rect 40271 32388 40316 32416
rect 40129 32379 40187 32385
rect 40310 32376 40316 32388
rect 40368 32376 40374 32428
rect 40972 32425 41000 32456
rect 40773 32419 40831 32425
rect 40773 32385 40785 32419
rect 40819 32385 40831 32419
rect 40773 32379 40831 32385
rect 40957 32419 41015 32425
rect 40957 32385 40969 32419
rect 41003 32385 41015 32419
rect 40957 32379 41015 32385
rect 41601 32419 41659 32425
rect 41601 32385 41613 32419
rect 41647 32416 41659 32419
rect 41690 32416 41696 32428
rect 41647 32388 41696 32416
rect 41647 32385 41659 32388
rect 41601 32379 41659 32385
rect 40788 32348 40816 32379
rect 41690 32376 41696 32388
rect 41748 32376 41754 32428
rect 42426 32416 42432 32428
rect 42387 32388 42432 32416
rect 42426 32376 42432 32388
rect 42484 32376 42490 32428
rect 43530 32416 43536 32428
rect 43491 32388 43536 32416
rect 43530 32376 43536 32388
rect 43588 32376 43594 32428
rect 44361 32419 44419 32425
rect 44361 32385 44373 32419
rect 44407 32416 44419 32419
rect 44450 32416 44456 32428
rect 44407 32388 44456 32416
rect 44407 32385 44419 32388
rect 44361 32379 44419 32385
rect 44450 32376 44456 32388
rect 44508 32376 44514 32428
rect 47762 32416 47768 32428
rect 47723 32388 47768 32416
rect 47762 32376 47768 32388
rect 47820 32376 47826 32428
rect 38795 32320 40816 32348
rect 42521 32351 42579 32357
rect 38795 32317 38807 32320
rect 38749 32311 38807 32317
rect 42521 32317 42533 32351
rect 42567 32317 42579 32351
rect 43346 32348 43352 32360
rect 43307 32320 43352 32348
rect 42521 32311 42579 32317
rect 36188 32252 38700 32280
rect 42536 32280 42564 32311
rect 43346 32308 43352 32320
rect 43404 32308 43410 32360
rect 46474 32280 46480 32292
rect 42536 32252 46480 32280
rect 24946 32172 24952 32224
rect 25004 32212 25010 32224
rect 25133 32215 25191 32221
rect 25133 32212 25145 32215
rect 25004 32184 25145 32212
rect 25004 32172 25010 32184
rect 25133 32181 25145 32184
rect 25179 32181 25191 32215
rect 25133 32175 25191 32181
rect 28626 32172 28632 32224
rect 28684 32212 28690 32224
rect 30929 32215 30987 32221
rect 30929 32212 30941 32215
rect 28684 32184 30941 32212
rect 28684 32172 28690 32184
rect 30929 32181 30941 32184
rect 30975 32212 30987 32215
rect 32582 32212 32588 32224
rect 30975 32184 32588 32212
rect 30975 32181 30987 32184
rect 30929 32175 30987 32181
rect 32582 32172 32588 32184
rect 32640 32212 32646 32224
rect 33870 32212 33876 32224
rect 32640 32184 33876 32212
rect 32640 32172 32646 32184
rect 33870 32172 33876 32184
rect 33928 32172 33934 32224
rect 36188 32221 36216 32252
rect 46474 32240 46480 32252
rect 46532 32240 46538 32292
rect 36173 32215 36231 32221
rect 36173 32181 36185 32215
rect 36219 32181 36231 32215
rect 44174 32212 44180 32224
rect 44135 32184 44180 32212
rect 36173 32175 36231 32181
rect 44174 32172 44180 32184
rect 44232 32172 44238 32224
rect 47578 32212 47584 32224
rect 47539 32184 47584 32212
rect 47578 32172 47584 32184
rect 47636 32172 47642 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 2498 32008 2504 32020
rect 2459 31980 2504 32008
rect 2498 31968 2504 31980
rect 2556 31968 2562 32020
rect 26050 32008 26056 32020
rect 26011 31980 26056 32008
rect 26050 31968 26056 31980
rect 26108 31968 26114 32020
rect 29546 31968 29552 32020
rect 29604 32008 29610 32020
rect 33229 32011 33287 32017
rect 29604 31980 30788 32008
rect 29604 31968 29610 31980
rect 29270 31900 29276 31952
rect 29328 31940 29334 31952
rect 30760 31949 30788 31980
rect 33229 31977 33241 32011
rect 33275 32008 33287 32011
rect 35434 32008 35440 32020
rect 33275 31980 35440 32008
rect 33275 31977 33287 31980
rect 33229 31971 33287 31977
rect 29825 31943 29883 31949
rect 29825 31940 29837 31943
rect 29328 31912 29837 31940
rect 29328 31900 29334 31912
rect 29825 31909 29837 31912
rect 29871 31909 29883 31943
rect 29825 31903 29883 31909
rect 30745 31943 30803 31949
rect 30745 31909 30757 31943
rect 30791 31909 30803 31943
rect 30745 31903 30803 31909
rect 24394 31832 24400 31884
rect 24452 31872 24458 31884
rect 24673 31875 24731 31881
rect 24673 31872 24685 31875
rect 24452 31844 24685 31872
rect 24452 31832 24458 31844
rect 24673 31841 24685 31844
rect 24719 31841 24731 31875
rect 27614 31872 27620 31884
rect 27575 31844 27620 31872
rect 24673 31835 24731 31841
rect 27614 31832 27620 31844
rect 27672 31832 27678 31884
rect 29178 31872 29184 31884
rect 28644 31844 29184 31872
rect 2409 31807 2467 31813
rect 2409 31773 2421 31807
rect 2455 31804 2467 31807
rect 8570 31804 8576 31816
rect 2455 31776 8576 31804
rect 2455 31773 2467 31776
rect 2409 31767 2467 31773
rect 8570 31764 8576 31776
rect 8628 31764 8634 31816
rect 24946 31813 24952 31816
rect 24940 31804 24952 31813
rect 24907 31776 24952 31804
rect 24940 31767 24952 31776
rect 24946 31764 24952 31767
rect 25004 31764 25010 31816
rect 27798 31804 27804 31816
rect 27759 31776 27804 31804
rect 27798 31764 27804 31776
rect 27856 31764 27862 31816
rect 28350 31764 28356 31816
rect 28408 31804 28414 31816
rect 28644 31813 28672 31844
rect 29178 31832 29184 31844
rect 29236 31832 29242 31884
rect 29546 31872 29552 31884
rect 29507 31844 29552 31872
rect 29546 31832 29552 31844
rect 29604 31832 29610 31884
rect 28445 31807 28503 31813
rect 28445 31804 28457 31807
rect 28408 31776 28457 31804
rect 28408 31764 28414 31776
rect 28445 31773 28457 31776
rect 28491 31773 28503 31807
rect 28445 31767 28503 31773
rect 28629 31807 28687 31813
rect 28629 31773 28641 31807
rect 28675 31773 28687 31807
rect 28629 31767 28687 31773
rect 28905 31807 28963 31813
rect 28905 31773 28917 31807
rect 28951 31804 28963 31807
rect 28994 31804 29000 31816
rect 28951 31776 29000 31804
rect 28951 31773 28963 31776
rect 28905 31767 28963 31773
rect 28994 31764 29000 31776
rect 29052 31804 29058 31816
rect 29730 31804 29736 31816
rect 29052 31776 29736 31804
rect 29052 31764 29058 31776
rect 29730 31764 29736 31776
rect 29788 31764 29794 31816
rect 29840 31804 29868 31903
rect 30098 31832 30104 31884
rect 30156 31872 30162 31884
rect 30929 31875 30987 31881
rect 30929 31872 30941 31875
rect 30156 31844 30941 31872
rect 30156 31832 30162 31844
rect 30929 31841 30941 31844
rect 30975 31841 30987 31875
rect 33042 31872 33048 31884
rect 30929 31835 30987 31841
rect 32324 31844 33048 31872
rect 30469 31807 30527 31813
rect 30469 31804 30481 31807
rect 29840 31776 30481 31804
rect 30469 31773 30481 31776
rect 30515 31773 30527 31807
rect 30469 31767 30527 31773
rect 31294 31764 31300 31816
rect 31352 31804 31358 31816
rect 32324 31813 32352 31844
rect 33042 31832 33048 31844
rect 33100 31872 33106 31884
rect 33244 31872 33272 31971
rect 35434 31968 35440 31980
rect 35492 31968 35498 32020
rect 36170 32008 36176 32020
rect 36131 31980 36176 32008
rect 36170 31968 36176 31980
rect 36228 31968 36234 32020
rect 36630 31968 36636 32020
rect 36688 32008 36694 32020
rect 37553 32011 37611 32017
rect 37553 32008 37565 32011
rect 36688 31980 37565 32008
rect 36688 31968 36694 31980
rect 37553 31977 37565 31980
rect 37599 31977 37611 32011
rect 42794 32008 42800 32020
rect 42707 31980 42800 32008
rect 37553 31971 37611 31977
rect 42794 31968 42800 31980
rect 42852 32008 42858 32020
rect 43530 32008 43536 32020
rect 42852 31980 43536 32008
rect 42852 31968 42858 31980
rect 43530 31968 43536 31980
rect 43588 31968 43594 32020
rect 33778 31940 33784 31952
rect 33739 31912 33784 31940
rect 33778 31900 33784 31912
rect 33836 31900 33842 31952
rect 37274 31940 37280 31952
rect 35820 31912 37280 31940
rect 34698 31872 34704 31884
rect 33100 31844 33272 31872
rect 33796 31844 34704 31872
rect 33100 31832 33106 31844
rect 32217 31807 32275 31813
rect 32217 31804 32229 31807
rect 31352 31776 32229 31804
rect 31352 31764 31358 31776
rect 32217 31773 32229 31776
rect 32263 31773 32275 31807
rect 32217 31767 32275 31773
rect 32309 31807 32367 31813
rect 32309 31773 32321 31807
rect 32355 31773 32367 31807
rect 32309 31767 32367 31773
rect 28810 31736 28816 31748
rect 28723 31708 28816 31736
rect 28810 31696 28816 31708
rect 28868 31736 28874 31748
rect 30098 31736 30104 31748
rect 28868 31708 30104 31736
rect 28868 31696 28874 31708
rect 30098 31696 30104 31708
rect 30156 31696 30162 31748
rect 32232 31736 32260 31767
rect 32398 31764 32404 31816
rect 32456 31804 32462 31816
rect 32456 31776 32501 31804
rect 32456 31764 32462 31776
rect 32582 31764 32588 31816
rect 32640 31804 32646 31816
rect 32640 31776 32685 31804
rect 32640 31764 32646 31776
rect 32950 31764 32956 31816
rect 33008 31804 33014 31816
rect 33134 31804 33140 31816
rect 33008 31776 33140 31804
rect 33008 31764 33014 31776
rect 33134 31764 33140 31776
rect 33192 31764 33198 31816
rect 33796 31813 33824 31844
rect 34698 31832 34704 31844
rect 34756 31832 34762 31884
rect 33781 31807 33839 31813
rect 33781 31773 33793 31807
rect 33827 31773 33839 31807
rect 33781 31767 33839 31773
rect 34057 31807 34115 31813
rect 34057 31773 34069 31807
rect 34103 31804 34115 31807
rect 34422 31804 34428 31816
rect 34103 31776 34428 31804
rect 34103 31773 34115 31776
rect 34057 31767 34115 31773
rect 34422 31764 34428 31776
rect 34480 31804 34486 31816
rect 35820 31813 35848 31912
rect 37274 31900 37280 31912
rect 37332 31940 37338 31952
rect 37642 31940 37648 31952
rect 37332 31912 37648 31940
rect 37332 31900 37338 31912
rect 37642 31900 37648 31912
rect 37700 31940 37706 31952
rect 37921 31943 37979 31949
rect 37921 31940 37933 31943
rect 37700 31912 37933 31940
rect 37700 31900 37706 31912
rect 37921 31909 37933 31912
rect 37967 31909 37979 31943
rect 37921 31903 37979 31909
rect 38378 31900 38384 31952
rect 38436 31940 38442 31952
rect 42153 31943 42211 31949
rect 38436 31912 38700 31940
rect 38436 31900 38442 31912
rect 35894 31832 35900 31884
rect 35952 31872 35958 31884
rect 35952 31844 35997 31872
rect 35952 31832 35958 31844
rect 36998 31832 37004 31884
rect 37056 31872 37062 31884
rect 38010 31872 38016 31884
rect 37056 31844 37596 31872
rect 37971 31844 38016 31872
rect 37056 31832 37062 31844
rect 35805 31807 35863 31813
rect 34480 31776 35572 31804
rect 34480 31764 34486 31776
rect 34146 31736 34152 31748
rect 32232 31708 34152 31736
rect 34146 31696 34152 31708
rect 34204 31696 34210 31748
rect 35544 31736 35572 31776
rect 35805 31773 35817 31807
rect 35851 31773 35863 31807
rect 35805 31767 35863 31773
rect 36538 31764 36544 31816
rect 36596 31804 36602 31816
rect 36633 31807 36691 31813
rect 36633 31804 36645 31807
rect 36596 31776 36645 31804
rect 36596 31764 36602 31776
rect 36633 31773 36645 31776
rect 36679 31773 36691 31807
rect 36633 31767 36691 31773
rect 36817 31807 36875 31813
rect 36817 31773 36829 31807
rect 36863 31782 36875 31807
rect 37090 31804 37096 31816
rect 36906 31782 36912 31794
rect 36863 31773 36912 31782
rect 36817 31767 36912 31773
rect 36832 31754 36912 31767
rect 36832 31736 36860 31754
rect 36906 31742 36912 31754
rect 36964 31742 36970 31794
rect 37051 31776 37096 31804
rect 37090 31764 37096 31776
rect 37148 31764 37154 31816
rect 37568 31770 37596 31844
rect 38010 31832 38016 31844
rect 38068 31832 38074 31884
rect 37737 31807 37795 31813
rect 37737 31773 37749 31807
rect 37783 31804 37795 31807
rect 38562 31804 38568 31816
rect 37783 31776 38568 31804
rect 37783 31773 37795 31776
rect 37568 31742 37688 31770
rect 37737 31767 37795 31773
rect 38562 31764 38568 31776
rect 38620 31764 38626 31816
rect 38672 31745 38700 31912
rect 42153 31909 42165 31943
rect 42199 31940 42211 31943
rect 42518 31940 42524 31952
rect 42199 31912 42524 31940
rect 42199 31909 42211 31912
rect 42153 31903 42211 31909
rect 42518 31900 42524 31912
rect 42576 31900 42582 31952
rect 46934 31940 46940 31952
rect 46308 31912 46940 31940
rect 39942 31872 39948 31884
rect 39903 31844 39948 31872
rect 39942 31832 39948 31844
rect 40000 31832 40006 31884
rect 40402 31872 40408 31884
rect 40363 31844 40408 31872
rect 40402 31832 40408 31844
rect 40460 31832 40466 31884
rect 41690 31832 41696 31884
rect 41748 31872 41754 31884
rect 41748 31844 43024 31872
rect 41748 31832 41754 31844
rect 40034 31804 40040 31816
rect 39995 31776 40040 31804
rect 40034 31764 40040 31776
rect 40092 31764 40098 31816
rect 41414 31764 41420 31816
rect 41472 31804 41478 31816
rect 42334 31804 42340 31816
rect 41472 31776 41517 31804
rect 42295 31776 42340 31804
rect 41472 31764 41478 31776
rect 42334 31764 42340 31776
rect 42392 31764 42398 31816
rect 42996 31813 43024 31844
rect 42981 31807 43039 31813
rect 42981 31773 42993 31807
rect 43027 31804 43039 31807
rect 43438 31804 43444 31816
rect 43027 31776 43444 31804
rect 43027 31773 43039 31776
rect 42981 31767 43039 31773
rect 43438 31764 43444 31776
rect 43496 31764 43502 31816
rect 46308 31813 46336 31912
rect 46934 31900 46940 31912
rect 46992 31900 46998 31952
rect 46474 31872 46480 31884
rect 46435 31844 46480 31872
rect 46474 31832 46480 31844
rect 46532 31832 46538 31884
rect 48130 31872 48136 31884
rect 48091 31844 48136 31872
rect 48130 31832 48136 31844
rect 48188 31832 48194 31884
rect 46293 31807 46351 31813
rect 46293 31773 46305 31807
rect 46339 31773 46351 31807
rect 46293 31767 46351 31773
rect 35544 31708 36860 31736
rect 37660 31736 37688 31742
rect 38473 31739 38531 31745
rect 38473 31736 38485 31739
rect 37660 31708 38485 31736
rect 38473 31705 38485 31708
rect 38519 31705 38531 31739
rect 38473 31699 38531 31705
rect 38657 31739 38715 31745
rect 38657 31705 38669 31739
rect 38703 31736 38715 31739
rect 40310 31736 40316 31748
rect 38703 31708 40316 31736
rect 38703 31705 38715 31708
rect 38657 31699 38715 31705
rect 40310 31696 40316 31708
rect 40368 31696 40374 31748
rect 43622 31736 43628 31748
rect 43583 31708 43628 31736
rect 43622 31696 43628 31708
rect 43680 31696 43686 31748
rect 43809 31739 43867 31745
rect 43809 31736 43821 31739
rect 43732 31708 43821 31736
rect 27982 31668 27988 31680
rect 27943 31640 27988 31668
rect 27982 31628 27988 31640
rect 28040 31628 28046 31680
rect 28902 31628 28908 31680
rect 28960 31668 28966 31680
rect 30009 31671 30067 31677
rect 30009 31668 30021 31671
rect 28960 31640 30021 31668
rect 28960 31628 28966 31640
rect 30009 31637 30021 31640
rect 30055 31637 30067 31671
rect 30009 31631 30067 31637
rect 31941 31671 31999 31677
rect 31941 31637 31953 31671
rect 31987 31668 31999 31671
rect 32214 31668 32220 31680
rect 31987 31640 32220 31668
rect 31987 31637 31999 31640
rect 31941 31631 31999 31637
rect 32214 31628 32220 31640
rect 32272 31628 32278 31680
rect 33962 31668 33968 31680
rect 33923 31640 33968 31668
rect 33962 31628 33968 31640
rect 34020 31628 34026 31680
rect 36998 31668 37004 31680
rect 36959 31640 37004 31668
rect 36998 31628 37004 31640
rect 37056 31628 37062 31680
rect 38838 31668 38844 31680
rect 38799 31640 38844 31668
rect 38838 31628 38844 31640
rect 38896 31628 38902 31680
rect 41230 31668 41236 31680
rect 41191 31640 41236 31668
rect 41230 31628 41236 31640
rect 41288 31628 41294 31680
rect 43162 31628 43168 31680
rect 43220 31668 43226 31680
rect 43732 31668 43760 31708
rect 43809 31705 43821 31708
rect 43855 31705 43867 31739
rect 43809 31699 43867 31705
rect 43898 31668 43904 31680
rect 43220 31640 43760 31668
rect 43859 31640 43904 31668
rect 43220 31628 43226 31640
rect 43898 31628 43904 31640
rect 43956 31628 43962 31680
rect 43990 31628 43996 31680
rect 44048 31668 44054 31680
rect 44177 31671 44235 31677
rect 44048 31640 44093 31668
rect 44048 31628 44054 31640
rect 44177 31637 44189 31671
rect 44223 31668 44235 31671
rect 44266 31668 44272 31680
rect 44223 31640 44272 31668
rect 44223 31637 44235 31640
rect 44177 31631 44235 31637
rect 44266 31628 44272 31640
rect 44324 31628 44330 31680
rect 46934 31628 46940 31680
rect 46992 31668 46998 31680
rect 48038 31668 48044 31680
rect 46992 31640 48044 31668
rect 46992 31628 46998 31640
rect 48038 31628 48044 31640
rect 48096 31628 48102 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 26421 31467 26479 31473
rect 26421 31433 26433 31467
rect 26467 31464 26479 31467
rect 26467 31436 34744 31464
rect 26467 31433 26479 31436
rect 26421 31427 26479 31433
rect 33778 31405 33784 31408
rect 33772 31396 33784 31405
rect 28644 31368 30420 31396
rect 33739 31368 33784 31396
rect 23842 31328 23848 31340
rect 23803 31300 23848 31328
rect 23842 31288 23848 31300
rect 23900 31288 23906 31340
rect 24029 31331 24087 31337
rect 24029 31297 24041 31331
rect 24075 31328 24087 31331
rect 24210 31328 24216 31340
rect 24075 31300 24216 31328
rect 24075 31297 24087 31300
rect 24029 31291 24087 31297
rect 24210 31288 24216 31300
rect 24268 31288 24274 31340
rect 24394 31288 24400 31340
rect 24452 31328 24458 31340
rect 25041 31331 25099 31337
rect 25041 31328 25053 31331
rect 24452 31300 25053 31328
rect 24452 31288 24458 31300
rect 25041 31297 25053 31300
rect 25087 31297 25099 31331
rect 25041 31291 25099 31297
rect 25130 31288 25136 31340
rect 25188 31328 25194 31340
rect 28644 31337 28672 31368
rect 25297 31331 25355 31337
rect 25297 31328 25309 31331
rect 25188 31300 25309 31328
rect 25188 31288 25194 31300
rect 25297 31297 25309 31300
rect 25343 31297 25355 31331
rect 25297 31291 25355 31297
rect 28629 31331 28687 31337
rect 28629 31297 28641 31331
rect 28675 31297 28687 31331
rect 28629 31291 28687 31297
rect 28813 31331 28871 31337
rect 28813 31297 28825 31331
rect 28859 31328 28871 31331
rect 29086 31328 29092 31340
rect 28859 31300 29092 31328
rect 28859 31297 28871 31300
rect 28813 31291 28871 31297
rect 29086 31288 29092 31300
rect 29144 31288 29150 31340
rect 29181 31331 29239 31337
rect 29181 31297 29193 31331
rect 29227 31297 29239 31331
rect 29181 31291 29239 31297
rect 28902 31260 28908 31272
rect 28863 31232 28908 31260
rect 28902 31220 28908 31232
rect 28960 31220 28966 31272
rect 28997 31263 29055 31269
rect 28997 31229 29009 31263
rect 29043 31229 29055 31263
rect 29196 31260 29224 31291
rect 29730 31288 29736 31340
rect 29788 31328 29794 31340
rect 30009 31331 30067 31337
rect 30009 31328 30021 31331
rect 29788 31300 30021 31328
rect 29788 31288 29794 31300
rect 30009 31297 30021 31300
rect 30055 31297 30067 31331
rect 30009 31291 30067 31297
rect 30098 31288 30104 31340
rect 30156 31328 30162 31340
rect 30282 31328 30288 31340
rect 30156 31300 30201 31328
rect 30243 31300 30288 31328
rect 30156 31288 30162 31300
rect 30282 31288 30288 31300
rect 30340 31288 30346 31340
rect 30392 31337 30420 31368
rect 33772 31359 33784 31368
rect 33778 31356 33784 31359
rect 33836 31356 33842 31408
rect 30377 31331 30435 31337
rect 30377 31297 30389 31331
rect 30423 31297 30435 31331
rect 30377 31291 30435 31297
rect 30116 31260 30144 31288
rect 29196 31232 30144 31260
rect 30392 31260 30420 31291
rect 31754 31288 31760 31340
rect 31812 31328 31818 31340
rect 33505 31331 33563 31337
rect 33505 31328 33517 31331
rect 31812 31300 33517 31328
rect 31812 31288 31818 31300
rect 33505 31297 33517 31300
rect 33551 31297 33563 31331
rect 33505 31291 33563 31297
rect 32030 31260 32036 31272
rect 30392 31232 32036 31260
rect 28997 31223 29055 31229
rect 27982 31152 27988 31204
rect 28040 31192 28046 31204
rect 28442 31192 28448 31204
rect 28040 31164 28448 31192
rect 28040 31152 28046 31164
rect 28442 31152 28448 31164
rect 28500 31192 28506 31204
rect 29012 31192 29040 31223
rect 32030 31220 32036 31232
rect 32088 31220 32094 31272
rect 34716 31260 34744 31436
rect 34790 31424 34796 31476
rect 34848 31464 34854 31476
rect 34885 31467 34943 31473
rect 34885 31464 34897 31467
rect 34848 31436 34897 31464
rect 34848 31424 34854 31436
rect 34885 31433 34897 31436
rect 34931 31433 34943 31467
rect 34885 31427 34943 31433
rect 36725 31467 36783 31473
rect 36725 31433 36737 31467
rect 36771 31464 36783 31467
rect 36998 31464 37004 31476
rect 36771 31436 37004 31464
rect 36771 31433 36783 31436
rect 36725 31427 36783 31433
rect 36998 31424 37004 31436
rect 37056 31424 37062 31476
rect 42886 31424 42892 31476
rect 42944 31464 42950 31476
rect 43346 31464 43352 31476
rect 42944 31436 43352 31464
rect 42944 31424 42950 31436
rect 43346 31424 43352 31436
rect 43404 31464 43410 31476
rect 43990 31464 43996 31476
rect 43404 31436 43996 31464
rect 43404 31424 43410 31436
rect 43990 31424 43996 31436
rect 44048 31464 44054 31476
rect 45189 31467 45247 31473
rect 45189 31464 45201 31467
rect 44048 31436 45201 31464
rect 44048 31424 44054 31436
rect 45189 31433 45201 31436
rect 45235 31433 45247 31467
rect 46845 31467 46903 31473
rect 46845 31464 46857 31467
rect 45189 31427 45247 31433
rect 45756 31436 46857 31464
rect 36170 31356 36176 31408
rect 36228 31396 36234 31408
rect 36357 31399 36415 31405
rect 36357 31396 36369 31399
rect 36228 31368 36369 31396
rect 36228 31356 36234 31368
rect 36357 31365 36369 31368
rect 36403 31365 36415 31399
rect 36357 31359 36415 31365
rect 36446 31356 36452 31408
rect 36504 31396 36510 31408
rect 36541 31399 36599 31405
rect 36541 31396 36553 31399
rect 36504 31368 36553 31396
rect 36504 31356 36510 31368
rect 36541 31365 36553 31368
rect 36587 31365 36599 31399
rect 40402 31396 40408 31408
rect 36541 31359 36599 31365
rect 38764 31368 40408 31396
rect 36906 31288 36912 31340
rect 36964 31328 36970 31340
rect 38764 31337 38792 31368
rect 40402 31356 40408 31368
rect 40460 31356 40466 31408
rect 40764 31399 40822 31405
rect 40764 31365 40776 31399
rect 40810 31396 40822 31399
rect 41230 31396 41236 31408
rect 40810 31368 41236 31396
rect 40810 31365 40822 31368
rect 40764 31359 40822 31365
rect 41230 31356 41236 31368
rect 41288 31356 41294 31408
rect 43622 31396 43628 31408
rect 41386 31368 43628 31396
rect 38657 31331 38715 31337
rect 38657 31328 38669 31331
rect 36964 31300 38669 31328
rect 36964 31288 36970 31300
rect 38657 31297 38669 31300
rect 38703 31297 38715 31331
rect 38657 31291 38715 31297
rect 38749 31331 38807 31337
rect 38749 31297 38761 31331
rect 38795 31297 38807 31331
rect 38749 31291 38807 31297
rect 38838 31288 38844 31340
rect 38896 31328 38902 31340
rect 39022 31328 39028 31340
rect 38896 31300 38941 31328
rect 38983 31300 39028 31328
rect 38896 31288 38902 31300
rect 39022 31288 39028 31300
rect 39080 31288 39086 31340
rect 41138 31328 41144 31340
rect 39132 31300 41144 31328
rect 39132 31260 39160 31300
rect 41138 31288 41144 31300
rect 41196 31328 41202 31340
rect 41386 31328 41414 31368
rect 42886 31328 42892 31340
rect 41196 31300 41414 31328
rect 42847 31300 42892 31328
rect 41196 31288 41202 31300
rect 42886 31288 42892 31300
rect 42944 31288 42950 31340
rect 43180 31337 43208 31368
rect 43622 31356 43628 31368
rect 43680 31356 43686 31408
rect 44076 31399 44134 31405
rect 44076 31365 44088 31399
rect 44122 31396 44134 31399
rect 44174 31396 44180 31408
rect 44122 31368 44180 31396
rect 44122 31365 44134 31368
rect 44076 31359 44134 31365
rect 44174 31356 44180 31368
rect 44232 31356 44238 31408
rect 45756 31340 45784 31436
rect 46845 31433 46857 31436
rect 46891 31464 46903 31467
rect 47486 31464 47492 31476
rect 46891 31436 47492 31464
rect 46891 31433 46903 31436
rect 46845 31427 46903 31433
rect 47486 31424 47492 31436
rect 47544 31424 47550 31476
rect 47762 31424 47768 31476
rect 47820 31464 47826 31476
rect 47949 31467 48007 31473
rect 47949 31464 47961 31467
rect 47820 31436 47961 31464
rect 47820 31424 47826 31436
rect 47949 31433 47961 31436
rect 47995 31433 48007 31467
rect 47949 31427 48007 31433
rect 46106 31356 46112 31408
rect 46164 31396 46170 31408
rect 46477 31399 46535 31405
rect 46477 31396 46489 31399
rect 46164 31368 46489 31396
rect 46164 31356 46170 31368
rect 46477 31365 46489 31368
rect 46523 31365 46535 31399
rect 46477 31359 46535 31365
rect 46753 31399 46811 31405
rect 46753 31365 46765 31399
rect 46799 31396 46811 31399
rect 47026 31396 47032 31408
rect 46799 31368 47032 31396
rect 46799 31365 46811 31368
rect 46753 31359 46811 31365
rect 47026 31356 47032 31368
rect 47084 31356 47090 31408
rect 43165 31331 43223 31337
rect 43165 31297 43177 31331
rect 43211 31297 43223 31331
rect 43898 31328 43904 31340
rect 43165 31291 43223 31297
rect 43456 31300 43904 31328
rect 34716 31232 39160 31260
rect 40497 31263 40555 31269
rect 40497 31229 40509 31263
rect 40543 31229 40555 31263
rect 43070 31260 43076 31272
rect 42983 31232 43076 31260
rect 40497 31223 40555 31229
rect 28500 31164 29040 31192
rect 28500 31152 28506 31164
rect 38746 31152 38752 31204
rect 38804 31192 38810 31204
rect 40512 31192 40540 31223
rect 43070 31220 43076 31232
rect 43128 31260 43134 31272
rect 43456 31260 43484 31300
rect 43898 31288 43904 31300
rect 43956 31288 43962 31340
rect 45738 31328 45744 31340
rect 45651 31300 45744 31328
rect 45738 31288 45744 31300
rect 45796 31288 45802 31340
rect 45833 31331 45891 31337
rect 45833 31297 45845 31331
rect 45879 31297 45891 31331
rect 45833 31291 45891 31297
rect 43806 31260 43812 31272
rect 43128 31232 43484 31260
rect 43767 31232 43812 31260
rect 43128 31220 43134 31232
rect 43806 31220 43812 31232
rect 43864 31220 43870 31272
rect 45848 31260 45876 31291
rect 46014 31288 46020 31340
rect 46072 31328 46078 31340
rect 46661 31331 46719 31337
rect 46661 31328 46673 31331
rect 46072 31300 46673 31328
rect 46072 31288 46078 31300
rect 46661 31297 46673 31300
rect 46707 31328 46719 31331
rect 46842 31328 46848 31340
rect 46707 31300 46848 31328
rect 46707 31297 46719 31300
rect 46661 31291 46719 31297
rect 46842 31288 46848 31300
rect 46900 31288 46906 31340
rect 47302 31328 47308 31340
rect 47044 31300 47308 31328
rect 47044 31260 47072 31300
rect 47302 31288 47308 31300
rect 47360 31328 47366 31340
rect 47765 31331 47823 31337
rect 47765 31328 47777 31331
rect 47360 31300 47777 31328
rect 47360 31288 47366 31300
rect 47765 31297 47777 31300
rect 47811 31297 47823 31331
rect 47765 31291 47823 31297
rect 45848 31232 47072 31260
rect 47581 31263 47639 31269
rect 47581 31229 47593 31263
rect 47627 31260 47639 31263
rect 48038 31260 48044 31272
rect 47627 31232 48044 31260
rect 47627 31229 47639 31232
rect 47581 31223 47639 31229
rect 48038 31220 48044 31232
rect 48096 31220 48102 31272
rect 38804 31164 40540 31192
rect 38804 31152 38810 31164
rect 44818 31152 44824 31204
rect 44876 31192 44882 31204
rect 46017 31195 46075 31201
rect 44876 31164 45324 31192
rect 44876 31152 44882 31164
rect 24213 31127 24271 31133
rect 24213 31093 24225 31127
rect 24259 31124 24271 31127
rect 24854 31124 24860 31136
rect 24259 31096 24860 31124
rect 24259 31093 24271 31096
rect 24213 31087 24271 31093
rect 24854 31084 24860 31096
rect 24912 31084 24918 31136
rect 29270 31084 29276 31136
rect 29328 31124 29334 31136
rect 29365 31127 29423 31133
rect 29365 31124 29377 31127
rect 29328 31096 29377 31124
rect 29328 31084 29334 31096
rect 29365 31093 29377 31096
rect 29411 31093 29423 31127
rect 29822 31124 29828 31136
rect 29783 31096 29828 31124
rect 29365 31087 29423 31093
rect 29822 31084 29828 31096
rect 29880 31084 29886 31136
rect 33502 31084 33508 31136
rect 33560 31124 33566 31136
rect 34422 31124 34428 31136
rect 33560 31096 34428 31124
rect 33560 31084 33566 31096
rect 34422 31084 34428 31096
rect 34480 31084 34486 31136
rect 38381 31127 38439 31133
rect 38381 31093 38393 31127
rect 38427 31124 38439 31127
rect 38838 31124 38844 31136
rect 38427 31096 38844 31124
rect 38427 31093 38439 31096
rect 38381 31087 38439 31093
rect 38838 31084 38844 31096
rect 38896 31084 38902 31136
rect 41877 31127 41935 31133
rect 41877 31093 41889 31127
rect 41923 31124 41935 31127
rect 41966 31124 41972 31136
rect 41923 31096 41972 31124
rect 41923 31093 41935 31096
rect 41877 31087 41935 31093
rect 41966 31084 41972 31096
rect 42024 31124 42030 31136
rect 43162 31124 43168 31136
rect 42024 31096 43168 31124
rect 42024 31084 42030 31096
rect 43162 31084 43168 31096
rect 43220 31084 43226 31136
rect 43349 31127 43407 31133
rect 43349 31093 43361 31127
rect 43395 31124 43407 31127
rect 45094 31124 45100 31136
rect 43395 31096 45100 31124
rect 43395 31093 43407 31096
rect 43349 31087 43407 31093
rect 45094 31084 45100 31096
rect 45152 31084 45158 31136
rect 45296 31124 45324 31164
rect 46017 31161 46029 31195
rect 46063 31192 46075 31195
rect 47762 31192 47768 31204
rect 46063 31164 47768 31192
rect 46063 31161 46075 31164
rect 46017 31155 46075 31161
rect 47762 31152 47768 31164
rect 47820 31152 47826 31204
rect 47029 31127 47087 31133
rect 47029 31124 47041 31127
rect 45296 31096 47041 31124
rect 47029 31093 47041 31096
rect 47075 31093 47087 31127
rect 47029 31087 47087 31093
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 24673 30923 24731 30929
rect 24673 30889 24685 30923
rect 24719 30920 24731 30923
rect 25130 30920 25136 30932
rect 24719 30892 25136 30920
rect 24719 30889 24731 30892
rect 24673 30883 24731 30889
rect 25130 30880 25136 30892
rect 25188 30880 25194 30932
rect 28721 30923 28779 30929
rect 28721 30889 28733 30923
rect 28767 30920 28779 30923
rect 28902 30920 28908 30932
rect 28767 30892 28908 30920
rect 28767 30889 28779 30892
rect 28721 30883 28779 30889
rect 28902 30880 28908 30892
rect 28960 30880 28966 30932
rect 33962 30880 33968 30932
rect 34020 30920 34026 30932
rect 34057 30923 34115 30929
rect 34057 30920 34069 30923
rect 34020 30892 34069 30920
rect 34020 30880 34026 30892
rect 34057 30889 34069 30892
rect 34103 30889 34115 30923
rect 34698 30920 34704 30932
rect 34659 30892 34704 30920
rect 34057 30883 34115 30889
rect 34698 30880 34704 30892
rect 34756 30880 34762 30932
rect 41414 30880 41420 30932
rect 41472 30920 41478 30932
rect 41509 30923 41567 30929
rect 41509 30920 41521 30923
rect 41472 30892 41521 30920
rect 41472 30880 41478 30892
rect 41509 30889 41521 30892
rect 41555 30889 41567 30923
rect 42334 30920 42340 30932
rect 42295 30892 42340 30920
rect 41509 30883 41567 30889
rect 42334 30880 42340 30892
rect 42392 30880 42398 30932
rect 43349 30923 43407 30929
rect 43349 30889 43361 30923
rect 43395 30920 43407 30923
rect 44450 30920 44456 30932
rect 43395 30892 44456 30920
rect 43395 30889 43407 30892
rect 43349 30883 43407 30889
rect 44450 30880 44456 30892
rect 44508 30880 44514 30932
rect 46014 30920 46020 30932
rect 45975 30892 46020 30920
rect 46014 30880 46020 30892
rect 46072 30880 46078 30932
rect 47026 30920 47032 30932
rect 46124 30892 47032 30920
rect 43809 30855 43867 30861
rect 43809 30821 43821 30855
rect 43855 30852 43867 30855
rect 44174 30852 44180 30864
rect 43855 30824 44180 30852
rect 43855 30821 43867 30824
rect 43809 30815 43867 30821
rect 44174 30812 44180 30824
rect 44232 30812 44238 30864
rect 46124 30852 46152 30892
rect 47026 30880 47032 30892
rect 47084 30880 47090 30932
rect 47486 30880 47492 30932
rect 47544 30920 47550 30932
rect 48133 30923 48191 30929
rect 48133 30920 48145 30923
rect 47544 30892 48145 30920
rect 47544 30880 47550 30892
rect 48133 30889 48145 30892
rect 48179 30889 48191 30923
rect 48133 30883 48191 30889
rect 45940 30824 46152 30852
rect 33134 30744 33140 30796
rect 33192 30784 33198 30796
rect 39850 30784 39856 30796
rect 33192 30756 35204 30784
rect 33192 30744 33198 30756
rect 24854 30716 24860 30728
rect 24815 30688 24860 30716
rect 24854 30676 24860 30688
rect 24912 30676 24918 30728
rect 28442 30716 28448 30728
rect 28403 30688 28448 30716
rect 28442 30676 28448 30688
rect 28500 30676 28506 30728
rect 28537 30719 28595 30725
rect 28537 30685 28549 30719
rect 28583 30685 28595 30719
rect 28810 30716 28816 30728
rect 28771 30688 28816 30716
rect 28537 30679 28595 30685
rect 28552 30648 28580 30679
rect 28810 30676 28816 30688
rect 28868 30676 28874 30728
rect 32122 30716 32128 30728
rect 32083 30688 32128 30716
rect 32122 30676 32128 30688
rect 32180 30676 32186 30728
rect 32214 30676 32220 30728
rect 32272 30716 32278 30728
rect 32381 30719 32439 30725
rect 32381 30716 32393 30719
rect 32272 30688 32393 30716
rect 32272 30676 32278 30688
rect 32381 30685 32393 30688
rect 32427 30685 32439 30719
rect 32381 30679 32439 30685
rect 33965 30719 34023 30725
rect 33965 30685 33977 30719
rect 34011 30716 34023 30719
rect 34790 30716 34796 30728
rect 34011 30688 34796 30716
rect 34011 30685 34023 30688
rect 33965 30679 34023 30685
rect 34790 30676 34796 30688
rect 34848 30676 34854 30728
rect 35176 30725 35204 30756
rect 39040 30756 39856 30784
rect 34885 30719 34943 30725
rect 34885 30685 34897 30719
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 35161 30719 35219 30725
rect 35161 30685 35173 30719
rect 35207 30685 35219 30719
rect 35161 30679 35219 30685
rect 28994 30648 29000 30660
rect 28552 30620 29000 30648
rect 28994 30608 29000 30620
rect 29052 30608 29058 30660
rect 27430 30540 27436 30592
rect 27488 30580 27494 30592
rect 28261 30583 28319 30589
rect 28261 30580 28273 30583
rect 27488 30552 28273 30580
rect 27488 30540 27494 30552
rect 28261 30549 28273 30552
rect 28307 30549 28319 30583
rect 33502 30580 33508 30592
rect 33463 30552 33508 30580
rect 28261 30543 28319 30549
rect 33502 30540 33508 30552
rect 33560 30540 33566 30592
rect 34900 30580 34928 30679
rect 39040 30660 39068 30756
rect 39850 30744 39856 30756
rect 39908 30784 39914 30796
rect 41598 30784 41604 30796
rect 39908 30756 41604 30784
rect 39908 30744 39914 30756
rect 41598 30744 41604 30756
rect 41656 30744 41662 30796
rect 41966 30784 41972 30796
rect 41927 30756 41972 30784
rect 41966 30744 41972 30756
rect 42024 30744 42030 30796
rect 42794 30784 42800 30796
rect 42168 30756 42800 30784
rect 40126 30676 40132 30728
rect 40184 30716 40190 30728
rect 40313 30719 40371 30725
rect 40313 30716 40325 30719
rect 40184 30688 40325 30716
rect 40184 30676 40190 30688
rect 40313 30685 40325 30688
rect 40359 30685 40371 30719
rect 41138 30716 41144 30728
rect 41099 30688 41144 30716
rect 40313 30679 40371 30685
rect 41138 30676 41144 30688
rect 41196 30676 41202 30728
rect 41325 30719 41383 30725
rect 41325 30685 41337 30719
rect 41371 30716 41383 30719
rect 41414 30716 41420 30728
rect 41371 30688 41420 30716
rect 41371 30685 41383 30688
rect 41325 30679 41383 30685
rect 41414 30676 41420 30688
rect 41472 30716 41478 30728
rect 42168 30725 42196 30756
rect 42794 30744 42800 30756
rect 42852 30784 42858 30796
rect 44266 30784 44272 30796
rect 42852 30756 43208 30784
rect 42852 30744 42858 30756
rect 42153 30719 42211 30725
rect 42153 30716 42165 30719
rect 41472 30688 42165 30716
rect 41472 30676 41478 30688
rect 42153 30685 42165 30688
rect 42199 30685 42211 30719
rect 43070 30716 43076 30728
rect 43031 30688 43076 30716
rect 42153 30679 42211 30685
rect 43070 30676 43076 30688
rect 43128 30676 43134 30728
rect 43180 30725 43208 30756
rect 44008 30756 44272 30784
rect 44008 30725 44036 30756
rect 44266 30744 44272 30756
rect 44324 30744 44330 30796
rect 44358 30744 44364 30796
rect 44416 30744 44422 30796
rect 45940 30793 45968 30824
rect 45925 30787 45983 30793
rect 45925 30753 45937 30787
rect 45971 30753 45983 30787
rect 46753 30787 46811 30793
rect 46753 30784 46765 30787
rect 45925 30747 45983 30753
rect 46032 30756 46765 30784
rect 43165 30719 43223 30725
rect 43165 30685 43177 30719
rect 43211 30685 43223 30719
rect 43165 30679 43223 30685
rect 43993 30719 44051 30725
rect 43993 30685 44005 30719
rect 44039 30685 44051 30719
rect 43993 30679 44051 30685
rect 44177 30719 44235 30725
rect 44177 30685 44189 30719
rect 44223 30716 44235 30719
rect 44376 30716 44404 30744
rect 44223 30688 44404 30716
rect 44223 30685 44235 30688
rect 44177 30679 44235 30685
rect 44450 30676 44456 30728
rect 44508 30716 44514 30728
rect 45373 30719 45431 30725
rect 45373 30716 45385 30719
rect 44508 30688 44553 30716
rect 44836 30688 45385 30716
rect 44508 30676 44514 30688
rect 34974 30608 34980 30660
rect 35032 30648 35038 30660
rect 35069 30651 35127 30657
rect 35069 30648 35081 30651
rect 35032 30620 35081 30648
rect 35032 30608 35038 30620
rect 35069 30617 35081 30620
rect 35115 30617 35127 30651
rect 35069 30611 35127 30617
rect 36357 30651 36415 30657
rect 36357 30617 36369 30651
rect 36403 30648 36415 30651
rect 37182 30648 37188 30660
rect 36403 30620 37188 30648
rect 36403 30617 36415 30620
rect 36357 30611 36415 30617
rect 37182 30608 37188 30620
rect 37240 30608 37246 30660
rect 38102 30648 38108 30660
rect 38015 30620 38108 30648
rect 38102 30608 38108 30620
rect 38160 30648 38166 30660
rect 39022 30648 39028 30660
rect 38160 30620 39028 30648
rect 38160 30608 38166 30620
rect 39022 30608 39028 30620
rect 39080 30608 39086 30660
rect 44085 30651 44143 30657
rect 44085 30617 44097 30651
rect 44131 30617 44143 30651
rect 44085 30611 44143 30617
rect 44315 30651 44373 30657
rect 44315 30617 44327 30651
rect 44361 30648 44373 30651
rect 44836 30648 44864 30688
rect 45373 30685 45385 30688
rect 45419 30685 45431 30719
rect 45373 30679 45431 30685
rect 45646 30676 45652 30728
rect 45704 30716 45710 30728
rect 46032 30716 46060 30756
rect 46753 30753 46765 30756
rect 46799 30753 46811 30787
rect 46753 30747 46811 30753
rect 45704 30688 46060 30716
rect 45704 30676 45710 30688
rect 46106 30676 46112 30728
rect 46164 30716 46170 30728
rect 47020 30719 47078 30725
rect 46164 30688 46209 30716
rect 46164 30676 46170 30688
rect 47020 30685 47032 30719
rect 47066 30716 47078 30719
rect 47578 30716 47584 30728
rect 47066 30688 47584 30716
rect 47066 30685 47078 30688
rect 47020 30679 47078 30685
rect 47578 30676 47584 30688
rect 47636 30676 47642 30728
rect 44361 30620 44864 30648
rect 45005 30651 45063 30657
rect 44361 30617 44373 30620
rect 44315 30611 44373 30617
rect 45005 30617 45017 30651
rect 45051 30617 45063 30651
rect 45005 30611 45063 30617
rect 36262 30580 36268 30592
rect 34900 30552 36268 30580
rect 36262 30540 36268 30552
rect 36320 30540 36326 30592
rect 40402 30580 40408 30592
rect 40363 30552 40408 30580
rect 40402 30540 40408 30552
rect 40460 30580 40466 30592
rect 40586 30580 40592 30592
rect 40460 30552 40592 30580
rect 40460 30540 40466 30552
rect 40586 30540 40592 30552
rect 40644 30540 40650 30592
rect 44100 30580 44128 30611
rect 44818 30580 44824 30592
rect 44100 30552 44824 30580
rect 44818 30540 44824 30552
rect 44876 30540 44882 30592
rect 45020 30580 45048 30611
rect 45094 30608 45100 30660
rect 45152 30648 45158 30660
rect 45189 30651 45247 30657
rect 45189 30648 45201 30651
rect 45152 30620 45201 30648
rect 45152 30608 45158 30620
rect 45189 30617 45201 30620
rect 45235 30617 45247 30651
rect 45189 30611 45247 30617
rect 45738 30608 45744 30660
rect 45796 30648 45802 30660
rect 45833 30651 45891 30657
rect 45833 30648 45845 30651
rect 45796 30620 45845 30648
rect 45796 30608 45802 30620
rect 45833 30617 45845 30620
rect 45879 30617 45891 30651
rect 45833 30611 45891 30617
rect 46293 30583 46351 30589
rect 46293 30580 46305 30583
rect 45020 30552 46305 30580
rect 46293 30549 46305 30552
rect 46339 30549 46351 30583
rect 46293 30543 46351 30549
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 36004 30348 36584 30376
rect 30834 30268 30840 30320
rect 30892 30308 30898 30320
rect 31113 30311 31171 30317
rect 31113 30308 31125 30311
rect 30892 30280 31125 30308
rect 30892 30268 30898 30280
rect 31113 30277 31125 30280
rect 31159 30308 31171 30311
rect 36004 30308 36032 30348
rect 36556 30308 36584 30348
rect 38930 30336 38936 30388
rect 38988 30376 38994 30388
rect 41598 30376 41604 30388
rect 38988 30348 41604 30376
rect 38988 30336 38994 30348
rect 41598 30336 41604 30348
rect 41656 30336 41662 30388
rect 47026 30376 47032 30388
rect 46987 30348 47032 30376
rect 47026 30336 47032 30348
rect 47084 30336 47090 30388
rect 40402 30308 40408 30320
rect 31159 30280 36032 30308
rect 36280 30280 36492 30308
rect 36556 30280 40408 30308
rect 31159 30277 31171 30280
rect 31113 30271 31171 30277
rect 29270 30240 29276 30252
rect 29231 30212 29276 30240
rect 29270 30200 29276 30212
rect 29328 30200 29334 30252
rect 29454 30240 29460 30252
rect 29415 30212 29460 30240
rect 29454 30200 29460 30212
rect 29512 30200 29518 30252
rect 35434 30200 35440 30252
rect 35492 30240 35498 30252
rect 36280 30240 36308 30280
rect 36464 30249 36492 30280
rect 40402 30268 40408 30280
rect 40460 30268 40466 30320
rect 41414 30268 41420 30320
rect 41472 30308 41478 30320
rect 43806 30308 43812 30320
rect 41472 30280 41517 30308
rect 42444 30280 43812 30308
rect 41472 30268 41478 30280
rect 35492 30212 36308 30240
rect 36357 30243 36415 30249
rect 35492 30200 35498 30212
rect 36357 30209 36369 30243
rect 36403 30209 36415 30243
rect 36357 30203 36415 30209
rect 36449 30243 36507 30249
rect 36449 30209 36461 30243
rect 36495 30209 36507 30243
rect 36449 30203 36507 30209
rect 36372 30172 36400 30203
rect 36538 30200 36544 30252
rect 36596 30240 36602 30252
rect 36596 30212 36641 30240
rect 36596 30200 36602 30212
rect 36722 30200 36728 30252
rect 36780 30240 36786 30252
rect 37274 30240 37280 30252
rect 36780 30212 36825 30240
rect 37235 30212 37280 30240
rect 36780 30200 36786 30212
rect 37274 30200 37280 30212
rect 37332 30200 37338 30252
rect 37366 30200 37372 30252
rect 37424 30240 37430 30252
rect 37461 30243 37519 30249
rect 37461 30240 37473 30243
rect 37424 30212 37473 30240
rect 37424 30200 37430 30212
rect 37461 30209 37473 30212
rect 37507 30209 37519 30243
rect 37461 30203 37519 30209
rect 37550 30200 37556 30252
rect 37608 30240 37614 30252
rect 37691 30243 37749 30249
rect 37608 30212 37653 30240
rect 37608 30200 37614 30212
rect 37691 30209 37703 30243
rect 37737 30240 37749 30243
rect 38562 30240 38568 30252
rect 37737 30212 38568 30240
rect 37737 30209 37749 30212
rect 37691 30203 37749 30209
rect 38562 30200 38568 30212
rect 38620 30200 38626 30252
rect 38746 30240 38752 30252
rect 38707 30212 38752 30240
rect 38746 30200 38752 30212
rect 38804 30200 38810 30252
rect 38838 30200 38844 30252
rect 38896 30240 38902 30252
rect 42444 30249 42472 30280
rect 43806 30268 43812 30280
rect 43864 30268 43870 30320
rect 39005 30243 39063 30249
rect 39005 30240 39017 30243
rect 38896 30212 39017 30240
rect 38896 30200 38902 30212
rect 39005 30209 39017 30212
rect 39051 30209 39063 30243
rect 39005 30203 39063 30209
rect 42429 30243 42487 30249
rect 42429 30209 42441 30243
rect 42475 30209 42487 30243
rect 42429 30203 42487 30209
rect 42518 30200 42524 30252
rect 42576 30240 42582 30252
rect 42685 30243 42743 30249
rect 42685 30240 42697 30243
rect 42576 30212 42697 30240
rect 42576 30200 42582 30212
rect 42685 30209 42697 30212
rect 42731 30209 42743 30243
rect 42685 30203 42743 30209
rect 45916 30243 45974 30249
rect 45916 30209 45928 30243
rect 45962 30240 45974 30243
rect 47762 30240 47768 30252
rect 45962 30212 47624 30240
rect 47723 30212 47768 30240
rect 45962 30209 45974 30212
rect 45916 30203 45974 30209
rect 37292 30172 37320 30200
rect 36372 30144 37320 30172
rect 31297 30107 31355 30113
rect 31297 30073 31309 30107
rect 31343 30104 31355 30107
rect 33410 30104 33416 30116
rect 31343 30076 33416 30104
rect 31343 30073 31355 30076
rect 31297 30067 31355 30073
rect 33410 30064 33416 30076
rect 33468 30064 33474 30116
rect 37292 30104 37320 30144
rect 43806 30132 43812 30184
rect 43864 30172 43870 30184
rect 45646 30172 45652 30184
rect 43864 30144 45652 30172
rect 43864 30132 43870 30144
rect 45646 30132 45652 30144
rect 45704 30132 45710 30184
rect 37642 30104 37648 30116
rect 37292 30076 37648 30104
rect 37642 30064 37648 30076
rect 37700 30064 37706 30116
rect 40129 30107 40187 30113
rect 40129 30073 40141 30107
rect 40175 30104 40187 30107
rect 40310 30104 40316 30116
rect 40175 30076 40316 30104
rect 40175 30073 40187 30076
rect 40129 30067 40187 30073
rect 40310 30064 40316 30076
rect 40368 30064 40374 30116
rect 41598 30104 41604 30116
rect 41559 30076 41604 30104
rect 41598 30064 41604 30076
rect 41656 30064 41662 30116
rect 47596 30113 47624 30212
rect 47762 30200 47768 30212
rect 47820 30200 47826 30252
rect 47581 30107 47639 30113
rect 47581 30073 47593 30107
rect 47627 30073 47639 30107
rect 47581 30067 47639 30073
rect 29273 30039 29331 30045
rect 29273 30005 29285 30039
rect 29319 30036 29331 30039
rect 30006 30036 30012 30048
rect 29319 30008 30012 30036
rect 29319 30005 29331 30008
rect 29273 29999 29331 30005
rect 30006 29996 30012 30008
rect 30064 29996 30070 30048
rect 36078 30036 36084 30048
rect 36039 30008 36084 30036
rect 36078 29996 36084 30008
rect 36136 29996 36142 30048
rect 37826 30036 37832 30048
rect 37787 30008 37832 30036
rect 37826 29996 37832 30008
rect 37884 29996 37890 30048
rect 43809 30039 43867 30045
rect 43809 30005 43821 30039
rect 43855 30036 43867 30039
rect 43898 30036 43904 30048
rect 43855 30008 43904 30036
rect 43855 30005 43867 30008
rect 43809 29999 43867 30005
rect 43898 29996 43904 30008
rect 43956 29996 43962 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 36814 29792 36820 29844
rect 36872 29832 36878 29844
rect 38930 29832 38936 29844
rect 36872 29804 38936 29832
rect 36872 29792 36878 29804
rect 38930 29792 38936 29804
rect 38988 29792 38994 29844
rect 40494 29832 40500 29844
rect 40455 29804 40500 29832
rect 40494 29792 40500 29804
rect 40552 29792 40558 29844
rect 43438 29832 43444 29844
rect 43399 29804 43444 29832
rect 43438 29792 43444 29804
rect 43496 29792 43502 29844
rect 34701 29767 34759 29773
rect 34701 29733 34713 29767
rect 34747 29764 34759 29767
rect 35894 29764 35900 29776
rect 34747 29736 35900 29764
rect 34747 29733 34759 29736
rect 34701 29727 34759 29733
rect 35894 29724 35900 29736
rect 35952 29724 35958 29776
rect 40310 29764 40316 29776
rect 38948 29736 40316 29764
rect 29270 29696 29276 29708
rect 25056 29668 25728 29696
rect 22646 29588 22652 29640
rect 22704 29628 22710 29640
rect 24670 29628 24676 29640
rect 22704 29600 24676 29628
rect 22704 29588 22710 29600
rect 24670 29588 24676 29600
rect 24728 29588 24734 29640
rect 24762 29628 24820 29634
rect 24762 29594 24774 29628
rect 24808 29594 24820 29628
rect 24762 29588 24820 29594
rect 24854 29588 24860 29640
rect 24912 29637 24918 29640
rect 25056 29637 25084 29668
rect 24912 29628 24920 29637
rect 25041 29631 25099 29637
rect 24912 29600 24957 29628
rect 24912 29591 24920 29600
rect 25041 29597 25053 29631
rect 25087 29597 25099 29631
rect 25590 29628 25596 29640
rect 25551 29600 25596 29628
rect 25041 29591 25099 29597
rect 24912 29588 24918 29591
rect 25590 29588 25596 29600
rect 25648 29588 25654 29640
rect 25700 29628 25728 29668
rect 28736 29668 29276 29696
rect 26326 29628 26332 29640
rect 25700 29600 26332 29628
rect 26326 29588 26332 29600
rect 26384 29588 26390 29640
rect 28736 29637 28764 29668
rect 29270 29656 29276 29668
rect 29328 29656 29334 29708
rect 30006 29696 30012 29708
rect 29967 29668 30012 29696
rect 30006 29656 30012 29668
rect 30064 29656 30070 29708
rect 32950 29656 32956 29708
rect 33008 29696 33014 29708
rect 36173 29699 36231 29705
rect 36173 29696 36185 29699
rect 33008 29668 36185 29696
rect 33008 29656 33014 29668
rect 36173 29665 36185 29668
rect 36219 29665 36231 29699
rect 36173 29659 36231 29665
rect 37550 29656 37556 29708
rect 37608 29696 37614 29708
rect 38010 29696 38016 29708
rect 37608 29668 38016 29696
rect 37608 29656 37614 29668
rect 38010 29656 38016 29668
rect 38068 29696 38074 29708
rect 38657 29699 38715 29705
rect 38657 29696 38669 29699
rect 38068 29668 38669 29696
rect 38068 29656 38074 29668
rect 38657 29665 38669 29668
rect 38703 29665 38715 29699
rect 38657 29659 38715 29665
rect 28721 29631 28779 29637
rect 28721 29597 28733 29631
rect 28767 29597 28779 29631
rect 28721 29591 28779 29597
rect 28997 29631 29055 29637
rect 28997 29597 29009 29631
rect 29043 29628 29055 29631
rect 29822 29628 29828 29640
rect 29043 29600 29828 29628
rect 29043 29597 29055 29600
rect 28997 29591 29055 29597
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 30101 29631 30159 29637
rect 30101 29597 30113 29631
rect 30147 29597 30159 29631
rect 30101 29591 30159 29597
rect 30929 29631 30987 29637
rect 30929 29597 30941 29631
rect 30975 29628 30987 29631
rect 32122 29628 32128 29640
rect 30975 29600 32128 29628
rect 30975 29597 30987 29600
rect 30929 29591 30987 29597
rect 24780 29504 24808 29588
rect 24394 29492 24400 29504
rect 24355 29464 24400 29492
rect 24394 29452 24400 29464
rect 24452 29452 24458 29504
rect 24762 29452 24768 29504
rect 24820 29452 24826 29504
rect 24854 29452 24860 29504
rect 24912 29492 24918 29504
rect 25608 29492 25636 29588
rect 25866 29569 25872 29572
rect 25860 29560 25872 29569
rect 25827 29532 25872 29560
rect 25860 29523 25872 29532
rect 25866 29520 25872 29523
rect 25924 29520 25930 29572
rect 28905 29563 28963 29569
rect 28905 29529 28917 29563
rect 28951 29560 28963 29563
rect 30116 29560 30144 29591
rect 32122 29588 32128 29600
rect 32180 29628 32186 29640
rect 32968 29628 32996 29656
rect 32180 29600 32996 29628
rect 33045 29631 33103 29637
rect 32180 29588 32186 29600
rect 33045 29597 33057 29631
rect 33091 29597 33103 29631
rect 33045 29591 33103 29597
rect 33137 29631 33195 29637
rect 33137 29597 33149 29631
rect 33183 29597 33195 29631
rect 33137 29591 33195 29597
rect 33229 29631 33287 29637
rect 33229 29597 33241 29631
rect 33275 29597 33287 29631
rect 33410 29628 33416 29640
rect 33323 29600 33416 29628
rect 33229 29591 33287 29597
rect 31196 29563 31254 29569
rect 28951 29532 31156 29560
rect 28951 29529 28963 29532
rect 28905 29523 28963 29529
rect 24912 29464 25636 29492
rect 24912 29452 24918 29464
rect 25958 29452 25964 29504
rect 26016 29492 26022 29504
rect 26973 29495 27031 29501
rect 26973 29492 26985 29495
rect 26016 29464 26985 29492
rect 26016 29452 26022 29464
rect 26973 29461 26985 29464
rect 27019 29461 27031 29495
rect 26973 29455 27031 29461
rect 28537 29495 28595 29501
rect 28537 29461 28549 29495
rect 28583 29492 28595 29495
rect 28810 29492 28816 29504
rect 28583 29464 28816 29492
rect 28583 29461 28595 29464
rect 28537 29455 28595 29461
rect 28810 29452 28816 29464
rect 28868 29452 28874 29504
rect 30469 29495 30527 29501
rect 30469 29461 30481 29495
rect 30515 29492 30527 29495
rect 30926 29492 30932 29504
rect 30515 29464 30932 29492
rect 30515 29461 30527 29464
rect 30469 29455 30527 29461
rect 30926 29452 30932 29464
rect 30984 29452 30990 29504
rect 31128 29492 31156 29532
rect 31196 29529 31208 29563
rect 31242 29560 31254 29563
rect 32769 29563 32827 29569
rect 32769 29560 32781 29563
rect 31242 29532 32781 29560
rect 31242 29529 31254 29532
rect 31196 29523 31254 29529
rect 32769 29529 32781 29532
rect 32815 29529 32827 29563
rect 33060 29560 33088 29591
rect 32769 29523 32827 29529
rect 32876 29532 33088 29560
rect 31478 29492 31484 29504
rect 31128 29464 31484 29492
rect 31478 29452 31484 29464
rect 31536 29452 31542 29504
rect 32122 29452 32128 29504
rect 32180 29492 32186 29504
rect 32309 29495 32367 29501
rect 32309 29492 32321 29495
rect 32180 29464 32321 29492
rect 32180 29452 32186 29464
rect 32309 29461 32321 29464
rect 32355 29492 32367 29495
rect 32876 29492 32904 29532
rect 33152 29504 33180 29591
rect 33244 29504 33272 29591
rect 33410 29588 33416 29600
rect 33468 29588 33474 29640
rect 33502 29588 33508 29640
rect 33560 29628 33566 29640
rect 33965 29631 34023 29637
rect 33965 29628 33977 29631
rect 33560 29600 33977 29628
rect 33560 29588 33566 29600
rect 33965 29597 33977 29600
rect 34011 29628 34023 29631
rect 34330 29628 34336 29640
rect 34011 29600 34336 29628
rect 34011 29597 34023 29600
rect 33965 29591 34023 29597
rect 34330 29588 34336 29600
rect 34388 29588 34394 29640
rect 34698 29588 34704 29640
rect 34756 29628 34762 29640
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34756 29600 34897 29628
rect 34756 29588 34762 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 35161 29631 35219 29637
rect 35161 29597 35173 29631
rect 35207 29628 35219 29631
rect 35342 29628 35348 29640
rect 35207 29600 35348 29628
rect 35207 29597 35219 29600
rect 35161 29591 35219 29597
rect 35342 29588 35348 29600
rect 35400 29588 35406 29640
rect 36078 29588 36084 29640
rect 36136 29628 36142 29640
rect 36429 29631 36487 29637
rect 36429 29628 36441 29631
rect 36136 29600 36441 29628
rect 36136 29588 36142 29600
rect 36429 29597 36441 29600
rect 36475 29597 36487 29631
rect 36429 29591 36487 29597
rect 37366 29588 37372 29640
rect 37424 29628 37430 29640
rect 38381 29631 38439 29637
rect 38381 29628 38393 29631
rect 37424 29600 38393 29628
rect 37424 29588 37430 29600
rect 38381 29597 38393 29600
rect 38427 29597 38439 29631
rect 38562 29628 38568 29640
rect 38523 29600 38568 29628
rect 38381 29591 38439 29597
rect 38562 29588 38568 29600
rect 38620 29588 38626 29640
rect 38948 29637 38976 29736
rect 39960 29637 39988 29736
rect 40310 29724 40316 29736
rect 40368 29724 40374 29776
rect 38749 29631 38807 29637
rect 38749 29597 38761 29631
rect 38795 29597 38807 29631
rect 38749 29591 38807 29597
rect 38933 29631 38991 29637
rect 38933 29597 38945 29631
rect 38979 29597 38991 29631
rect 38933 29591 38991 29597
rect 39117 29631 39175 29637
rect 39117 29597 39129 29631
rect 39163 29628 39175 29631
rect 39842 29631 39900 29637
rect 39842 29628 39854 29631
rect 39163 29600 39854 29628
rect 39163 29597 39175 29600
rect 39117 29591 39175 29597
rect 39842 29597 39854 29600
rect 39888 29597 39900 29631
rect 39960 29631 40031 29637
rect 39960 29600 39985 29631
rect 39842 29591 39900 29597
rect 39973 29597 39985 29600
rect 40019 29597 40031 29631
rect 39973 29591 40031 29597
rect 40359 29631 40417 29637
rect 40359 29597 40371 29631
rect 40405 29628 40417 29631
rect 41138 29628 41144 29640
rect 40405 29600 41144 29628
rect 40405 29597 40417 29600
rect 40359 29591 40417 29597
rect 33428 29560 33456 29588
rect 33778 29560 33784 29572
rect 33428 29532 33784 29560
rect 33778 29520 33784 29532
rect 33836 29520 33842 29572
rect 34146 29560 34152 29572
rect 34107 29532 34152 29560
rect 34146 29520 34152 29532
rect 34204 29520 34210 29572
rect 38764 29560 38792 29591
rect 41138 29588 41144 29600
rect 41196 29588 41202 29640
rect 43438 29588 43444 29640
rect 43496 29628 43502 29640
rect 44177 29631 44235 29637
rect 44177 29628 44189 29631
rect 43496 29600 44189 29628
rect 43496 29588 43502 29600
rect 44177 29597 44189 29600
rect 44223 29597 44235 29631
rect 46290 29628 46296 29640
rect 46251 29600 46296 29628
rect 44177 29591 44235 29597
rect 46290 29588 46296 29600
rect 46348 29588 46354 29640
rect 40126 29560 40132 29572
rect 38764 29532 40132 29560
rect 40126 29520 40132 29532
rect 40184 29520 40190 29572
rect 40218 29520 40224 29572
rect 40276 29560 40282 29572
rect 42613 29563 42671 29569
rect 40276 29532 40321 29560
rect 40276 29520 40282 29532
rect 42613 29529 42625 29563
rect 42659 29560 42671 29563
rect 43254 29560 43260 29572
rect 42659 29532 43260 29560
rect 42659 29529 42671 29532
rect 42613 29523 42671 29529
rect 43254 29520 43260 29532
rect 43312 29560 43318 29572
rect 43349 29563 43407 29569
rect 43349 29560 43361 29563
rect 43312 29532 43361 29560
rect 43312 29520 43318 29532
rect 43349 29529 43361 29532
rect 43395 29529 43407 29563
rect 46474 29560 46480 29572
rect 46435 29532 46480 29560
rect 43349 29523 43407 29529
rect 46474 29520 46480 29532
rect 46532 29520 46538 29572
rect 48130 29560 48136 29572
rect 48091 29532 48136 29560
rect 48130 29520 48136 29532
rect 48188 29520 48194 29572
rect 32355 29464 32904 29492
rect 32355 29461 32367 29464
rect 32309 29455 32367 29461
rect 33134 29452 33140 29504
rect 33192 29452 33198 29504
rect 33226 29452 33232 29504
rect 33284 29452 33290 29504
rect 33594 29452 33600 29504
rect 33652 29492 33658 29504
rect 35069 29495 35127 29501
rect 35069 29492 35081 29495
rect 33652 29464 35081 29492
rect 33652 29452 33658 29464
rect 35069 29461 35081 29464
rect 35115 29461 35127 29495
rect 35069 29455 35127 29461
rect 37274 29452 37280 29504
rect 37332 29492 37338 29504
rect 37553 29495 37611 29501
rect 37553 29492 37565 29495
rect 37332 29464 37565 29492
rect 37332 29452 37338 29464
rect 37553 29461 37565 29464
rect 37599 29461 37611 29495
rect 37553 29455 37611 29461
rect 37918 29452 37924 29504
rect 37976 29492 37982 29504
rect 42705 29495 42763 29501
rect 42705 29492 42717 29495
rect 37976 29464 42717 29492
rect 37976 29452 37982 29464
rect 42705 29461 42717 29464
rect 42751 29461 42763 29495
rect 42705 29455 42763 29461
rect 43993 29495 44051 29501
rect 43993 29461 44005 29495
rect 44039 29492 44051 29495
rect 44266 29492 44272 29504
rect 44039 29464 44272 29492
rect 44039 29461 44051 29464
rect 43993 29455 44051 29461
rect 44266 29452 44272 29464
rect 44324 29492 44330 29504
rect 44450 29492 44456 29504
rect 44324 29464 44456 29492
rect 44324 29452 44330 29464
rect 44450 29452 44456 29464
rect 44508 29452 44514 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 18874 29288 18880 29300
rect 18340 29260 18880 29288
rect 18340 29229 18368 29260
rect 18874 29248 18880 29260
rect 18932 29288 18938 29300
rect 24578 29288 24584 29300
rect 18932 29260 24584 29288
rect 18932 29248 18938 29260
rect 24578 29248 24584 29260
rect 24636 29248 24642 29300
rect 24670 29248 24676 29300
rect 24728 29288 24734 29300
rect 25225 29291 25283 29297
rect 25225 29288 25237 29291
rect 24728 29260 25237 29288
rect 24728 29248 24734 29260
rect 25225 29257 25237 29260
rect 25271 29257 25283 29291
rect 25225 29251 25283 29257
rect 25685 29291 25743 29297
rect 25685 29257 25697 29291
rect 25731 29288 25743 29291
rect 25866 29288 25872 29300
rect 25731 29260 25872 29288
rect 25731 29257 25743 29260
rect 25685 29251 25743 29257
rect 25866 29248 25872 29260
rect 25924 29248 25930 29300
rect 26234 29248 26240 29300
rect 26292 29248 26298 29300
rect 27614 29248 27620 29300
rect 27672 29288 27678 29300
rect 27672 29260 29408 29288
rect 27672 29248 27678 29260
rect 18325 29223 18383 29229
rect 18325 29189 18337 29223
rect 18371 29189 18383 29223
rect 24854 29220 24860 29232
rect 18325 29183 18383 29189
rect 23860 29192 24860 29220
rect 17770 29152 17776 29164
rect 17731 29124 17776 29152
rect 17770 29112 17776 29124
rect 17828 29112 17834 29164
rect 22833 29155 22891 29161
rect 22833 29121 22845 29155
rect 22879 29152 22891 29155
rect 23198 29152 23204 29164
rect 22879 29124 23204 29152
rect 22879 29121 22891 29124
rect 22833 29115 22891 29121
rect 23198 29112 23204 29124
rect 23256 29112 23262 29164
rect 23860 29161 23888 29192
rect 24854 29180 24860 29192
rect 24912 29180 24918 29232
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29121 23903 29155
rect 23845 29115 23903 29121
rect 24112 29155 24170 29161
rect 24112 29121 24124 29155
rect 24158 29152 24170 29155
rect 24394 29152 24400 29164
rect 24158 29124 24400 29152
rect 24158 29121 24170 29124
rect 24112 29115 24170 29121
rect 24394 29112 24400 29124
rect 24452 29112 24458 29164
rect 25866 29112 25872 29164
rect 25924 29161 25930 29164
rect 25924 29155 25973 29161
rect 25924 29121 25927 29155
rect 25961 29121 25973 29155
rect 25924 29115 25973 29121
rect 26066 29158 26124 29164
rect 26166 29158 26224 29161
rect 26252 29158 26280 29248
rect 29380 29220 29408 29260
rect 29454 29248 29460 29300
rect 29512 29288 29518 29300
rect 30009 29291 30067 29297
rect 30009 29288 30021 29291
rect 29512 29260 30021 29288
rect 29512 29248 29518 29260
rect 30009 29257 30021 29260
rect 30055 29257 30067 29291
rect 30009 29251 30067 29257
rect 31113 29291 31171 29297
rect 31113 29257 31125 29291
rect 31159 29288 31171 29291
rect 33226 29288 33232 29300
rect 31159 29260 33232 29288
rect 31159 29257 31171 29260
rect 31113 29251 31171 29257
rect 33226 29248 33232 29260
rect 33284 29248 33290 29300
rect 33321 29291 33379 29297
rect 33321 29257 33333 29291
rect 33367 29288 33379 29291
rect 35342 29288 35348 29300
rect 33367 29260 35020 29288
rect 35303 29260 35348 29288
rect 33367 29257 33379 29260
rect 33321 29251 33379 29257
rect 32122 29220 32128 29232
rect 29380 29192 30052 29220
rect 26066 29124 26078 29158
rect 26112 29124 26124 29158
rect 26160 29155 26280 29158
rect 26160 29124 26178 29155
rect 26066 29118 26124 29124
rect 26166 29121 26178 29124
rect 26212 29130 26280 29155
rect 26212 29121 26224 29130
rect 25924 29112 25930 29115
rect 22646 29084 22652 29096
rect 22607 29056 22652 29084
rect 22646 29044 22652 29056
rect 22704 29044 22710 29096
rect 25774 29044 25780 29096
rect 25832 29084 25838 29096
rect 26068 29084 26096 29118
rect 26166 29115 26224 29121
rect 26326 29112 26332 29164
rect 26384 29152 26390 29164
rect 27430 29152 27436 29164
rect 26384 29124 26477 29152
rect 27391 29124 27436 29152
rect 26384 29112 26390 29124
rect 27430 29112 27436 29124
rect 27488 29112 27494 29164
rect 28074 29152 28080 29164
rect 28035 29124 28080 29152
rect 28074 29112 28080 29124
rect 28132 29112 28138 29164
rect 28166 29112 28172 29164
rect 28224 29152 28230 29164
rect 28333 29155 28391 29161
rect 28333 29152 28345 29155
rect 28224 29124 28345 29152
rect 28224 29112 28230 29124
rect 28333 29121 28345 29124
rect 28379 29121 28391 29155
rect 29914 29152 29920 29164
rect 29875 29124 29920 29152
rect 28333 29115 28391 29121
rect 29914 29112 29920 29124
rect 29972 29112 29978 29164
rect 25832 29056 26096 29084
rect 26344 29084 26372 29112
rect 30024 29084 30052 29192
rect 30116 29192 32128 29220
rect 30116 29161 30144 29192
rect 32122 29180 32128 29192
rect 32180 29180 32186 29232
rect 33594 29180 33600 29232
rect 33652 29220 33658 29232
rect 33781 29223 33839 29229
rect 33781 29220 33793 29223
rect 33652 29192 33793 29220
rect 33652 29180 33658 29192
rect 33781 29189 33793 29192
rect 33827 29189 33839 29223
rect 34422 29220 34428 29232
rect 33781 29183 33839 29189
rect 34072 29192 34428 29220
rect 30101 29155 30159 29161
rect 30101 29121 30113 29155
rect 30147 29121 30159 29155
rect 30926 29152 30932 29164
rect 30887 29124 30932 29152
rect 30101 29115 30159 29121
rect 30926 29112 30932 29124
rect 30984 29112 30990 29164
rect 31113 29155 31171 29161
rect 31113 29121 31125 29155
rect 31159 29152 31171 29155
rect 31754 29152 31760 29164
rect 31159 29124 31760 29152
rect 31159 29121 31171 29124
rect 31113 29115 31171 29121
rect 31128 29084 31156 29115
rect 31754 29112 31760 29124
rect 31812 29112 31818 29164
rect 33137 29155 33195 29161
rect 33137 29121 33149 29155
rect 33183 29121 33195 29155
rect 33137 29115 33195 29121
rect 33321 29155 33379 29161
rect 33321 29121 33333 29155
rect 33367 29152 33379 29155
rect 33686 29152 33692 29164
rect 33367 29124 33692 29152
rect 33367 29121 33379 29124
rect 33321 29115 33379 29121
rect 26344 29056 27660 29084
rect 30024 29056 31156 29084
rect 33152 29084 33180 29115
rect 33686 29112 33692 29124
rect 33744 29112 33750 29164
rect 34072 29161 34100 29192
rect 34422 29180 34428 29192
rect 34480 29220 34486 29232
rect 34992 29229 35020 29260
rect 35342 29248 35348 29260
rect 35400 29248 35406 29300
rect 41138 29288 41144 29300
rect 41099 29260 41144 29288
rect 41138 29248 41144 29260
rect 41196 29248 41202 29300
rect 43438 29288 43444 29300
rect 43399 29260 43444 29288
rect 43438 29248 43444 29260
rect 43496 29248 43502 29300
rect 45002 29288 45008 29300
rect 44008 29260 45008 29288
rect 34977 29223 35035 29229
rect 34480 29192 34928 29220
rect 34480 29180 34486 29192
rect 34330 29161 34336 29164
rect 33965 29155 34023 29161
rect 33965 29121 33977 29155
rect 34011 29121 34023 29155
rect 33965 29115 34023 29121
rect 34057 29155 34115 29161
rect 34057 29121 34069 29155
rect 34103 29121 34115 29155
rect 34057 29115 34115 29121
rect 34315 29155 34336 29161
rect 34315 29121 34327 29155
rect 34315 29115 34336 29121
rect 33502 29084 33508 29096
rect 33152 29056 33508 29084
rect 25832 29044 25838 29056
rect 23017 29019 23075 29025
rect 23017 28985 23029 29019
rect 23063 29016 23075 29019
rect 23474 29016 23480 29028
rect 23063 28988 23480 29016
rect 23063 28985 23075 28988
rect 23017 28979 23075 28985
rect 23474 28976 23480 28988
rect 23532 28976 23538 29028
rect 26050 28976 26056 29028
rect 26108 29016 26114 29028
rect 26108 28988 26832 29016
rect 26108 28976 26114 28988
rect 22922 28908 22928 28960
rect 22980 28948 22986 28960
rect 26694 28948 26700 28960
rect 22980 28920 26700 28948
rect 22980 28908 22986 28920
rect 26694 28908 26700 28920
rect 26752 28908 26758 28960
rect 26804 28948 26832 28988
rect 27522 28948 27528 28960
rect 26804 28920 27528 28948
rect 27522 28908 27528 28920
rect 27580 28908 27586 28960
rect 27632 28948 27660 29056
rect 33502 29044 33508 29056
rect 33560 29044 33566 29096
rect 28718 28948 28724 28960
rect 27632 28920 28724 28948
rect 28718 28908 28724 28920
rect 28776 28908 28782 28960
rect 29454 28948 29460 28960
rect 29415 28920 29460 28948
rect 29454 28908 29460 28920
rect 29512 28908 29518 28960
rect 33980 28948 34008 29115
rect 34330 29112 34336 29115
rect 34388 29112 34394 29164
rect 34790 29152 34796 29164
rect 34751 29124 34796 29152
rect 34790 29112 34796 29124
rect 34848 29112 34854 29164
rect 34900 29152 34928 29192
rect 34977 29189 34989 29223
rect 35023 29189 35035 29223
rect 34977 29183 35035 29189
rect 35894 29180 35900 29232
rect 35952 29220 35958 29232
rect 36998 29220 37004 29232
rect 35952 29192 37004 29220
rect 35952 29180 35958 29192
rect 36998 29180 37004 29192
rect 37056 29180 37062 29232
rect 44008 29220 44036 29260
rect 45002 29248 45008 29260
rect 45060 29288 45066 29300
rect 45281 29291 45339 29297
rect 45281 29288 45293 29291
rect 45060 29260 45293 29288
rect 45060 29248 45066 29260
rect 45281 29257 45293 29260
rect 45327 29257 45339 29291
rect 45281 29251 45339 29257
rect 44174 29229 44180 29232
rect 44168 29220 44180 29229
rect 43180 29192 44036 29220
rect 44135 29192 44180 29220
rect 35069 29155 35127 29161
rect 35069 29152 35081 29155
rect 34900 29124 35081 29152
rect 35069 29121 35081 29124
rect 35115 29121 35127 29155
rect 35069 29115 35127 29121
rect 35161 29155 35219 29161
rect 35161 29121 35173 29155
rect 35207 29121 35219 29155
rect 36354 29152 36360 29164
rect 36315 29124 36360 29152
rect 35161 29115 35219 29121
rect 34422 29044 34428 29096
rect 34480 29084 34486 29096
rect 35176 29084 35204 29115
rect 36354 29112 36360 29124
rect 36412 29112 36418 29164
rect 36449 29155 36507 29161
rect 36449 29121 36461 29155
rect 36495 29121 36507 29155
rect 36449 29115 36507 29121
rect 36725 29155 36783 29161
rect 36725 29121 36737 29155
rect 36771 29152 36783 29155
rect 37274 29152 37280 29164
rect 36771 29124 37280 29152
rect 36771 29121 36783 29124
rect 36725 29115 36783 29121
rect 34480 29056 35204 29084
rect 34480 29044 34486 29056
rect 35986 29044 35992 29096
rect 36044 29084 36050 29096
rect 36464 29084 36492 29115
rect 37274 29112 37280 29124
rect 37332 29112 37338 29164
rect 37553 29155 37611 29161
rect 37553 29121 37565 29155
rect 37599 29152 37611 29155
rect 37642 29152 37648 29164
rect 37599 29124 37648 29152
rect 37599 29121 37611 29124
rect 37553 29115 37611 29121
rect 37642 29112 37648 29124
rect 37700 29112 37706 29164
rect 40129 29155 40187 29161
rect 40129 29121 40141 29155
rect 40175 29152 40187 29155
rect 40586 29152 40592 29164
rect 40175 29124 40592 29152
rect 40175 29121 40187 29124
rect 40129 29115 40187 29121
rect 40586 29112 40592 29124
rect 40644 29152 40650 29164
rect 43180 29161 43208 29192
rect 44168 29183 44180 29192
rect 44174 29180 44180 29183
rect 44232 29180 44238 29232
rect 41049 29155 41107 29161
rect 41049 29152 41061 29155
rect 40644 29124 41061 29152
rect 40644 29112 40650 29124
rect 41049 29121 41061 29124
rect 41095 29121 41107 29155
rect 41049 29115 41107 29121
rect 43165 29155 43223 29161
rect 43165 29121 43177 29155
rect 43211 29121 43223 29155
rect 43165 29115 43223 29121
rect 43257 29155 43315 29161
rect 43257 29121 43269 29155
rect 43303 29152 43315 29155
rect 43346 29152 43352 29164
rect 43303 29124 43352 29152
rect 43303 29121 43315 29124
rect 43257 29115 43315 29121
rect 43346 29112 43352 29124
rect 43404 29112 43410 29164
rect 46290 29112 46296 29164
rect 46348 29152 46354 29164
rect 47765 29155 47823 29161
rect 47765 29152 47777 29155
rect 46348 29124 47777 29152
rect 46348 29112 46354 29124
rect 47765 29121 47777 29124
rect 47811 29121 47823 29155
rect 47765 29115 47823 29121
rect 36044 29056 36492 29084
rect 36633 29087 36691 29093
rect 36044 29044 36050 29056
rect 36633 29053 36645 29087
rect 36679 29084 36691 29087
rect 37458 29084 37464 29096
rect 36679 29056 37464 29084
rect 36679 29053 36691 29056
rect 36633 29047 36691 29053
rect 37458 29044 37464 29056
rect 37516 29044 37522 29096
rect 43806 29044 43812 29096
rect 43864 29084 43870 29096
rect 43901 29087 43959 29093
rect 43901 29084 43913 29087
rect 43864 29056 43913 29084
rect 43864 29044 43870 29056
rect 43901 29053 43913 29056
rect 43947 29053 43959 29087
rect 43901 29047 43959 29053
rect 34238 28976 34244 29028
rect 34296 29016 34302 29028
rect 34296 28988 34341 29016
rect 34296 28976 34302 28988
rect 40494 28976 40500 29028
rect 40552 29016 40558 29028
rect 40589 29019 40647 29025
rect 40589 29016 40601 29019
rect 40552 28988 40601 29016
rect 40552 28976 40558 28988
rect 40589 28985 40601 28988
rect 40635 29016 40647 29019
rect 40770 29016 40776 29028
rect 40635 28988 40776 29016
rect 40635 28985 40647 28988
rect 40589 28979 40647 28985
rect 40770 28976 40776 28988
rect 40828 28976 40834 29028
rect 34422 28948 34428 28960
rect 33980 28920 34428 28948
rect 34422 28908 34428 28920
rect 34480 28908 34486 28960
rect 36170 28948 36176 28960
rect 36131 28920 36176 28948
rect 36170 28908 36176 28920
rect 36228 28908 36234 28960
rect 40218 28948 40224 28960
rect 40179 28920 40224 28948
rect 40218 28908 40224 28920
rect 40276 28908 40282 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 19978 28744 19984 28756
rect 19939 28716 19984 28744
rect 19978 28704 19984 28716
rect 20036 28704 20042 28756
rect 23753 28747 23811 28753
rect 23753 28713 23765 28747
rect 23799 28744 23811 28747
rect 24946 28744 24952 28756
rect 23799 28716 24952 28744
rect 23799 28713 23811 28716
rect 23753 28707 23811 28713
rect 24946 28704 24952 28716
rect 25004 28704 25010 28756
rect 26142 28704 26148 28756
rect 26200 28704 26206 28756
rect 26234 28704 26240 28756
rect 26292 28744 26298 28756
rect 26605 28747 26663 28753
rect 26605 28744 26617 28747
rect 26292 28716 26617 28744
rect 26292 28704 26298 28716
rect 26605 28713 26617 28716
rect 26651 28713 26663 28747
rect 26605 28707 26663 28713
rect 26694 28704 26700 28756
rect 26752 28744 26758 28756
rect 28077 28747 28135 28753
rect 26752 28716 27660 28744
rect 26752 28704 26758 28716
rect 23201 28679 23259 28685
rect 23201 28645 23213 28679
rect 23247 28645 23259 28679
rect 24762 28676 24768 28688
rect 24675 28648 24768 28676
rect 23201 28639 23259 28645
rect 18506 28608 18512 28620
rect 18467 28580 18512 28608
rect 18506 28568 18512 28580
rect 18564 28608 18570 28620
rect 18782 28608 18788 28620
rect 18564 28580 18788 28608
rect 18564 28568 18570 28580
rect 18782 28568 18788 28580
rect 18840 28568 18846 28620
rect 22925 28611 22983 28617
rect 22925 28577 22937 28611
rect 22971 28577 22983 28611
rect 22925 28571 22983 28577
rect 16853 28543 16911 28549
rect 16853 28509 16865 28543
rect 16899 28540 16911 28543
rect 22005 28543 22063 28549
rect 16899 28512 17816 28540
rect 16899 28509 16911 28512
rect 16853 28503 16911 28509
rect 17788 28484 17816 28512
rect 22005 28509 22017 28543
rect 22051 28540 22063 28543
rect 22646 28540 22652 28552
rect 22051 28512 22652 28540
rect 22051 28509 22063 28512
rect 22005 28503 22063 28509
rect 22646 28500 22652 28512
rect 22704 28500 22710 28552
rect 22830 28540 22836 28552
rect 22791 28512 22836 28540
rect 22830 28500 22836 28512
rect 22888 28500 22894 28552
rect 17126 28472 17132 28484
rect 17087 28444 17132 28472
rect 17126 28432 17132 28444
rect 17184 28432 17190 28484
rect 17770 28472 17776 28484
rect 17683 28444 17776 28472
rect 17770 28432 17776 28444
rect 17828 28472 17834 28484
rect 19705 28475 19763 28481
rect 19705 28472 19717 28475
rect 17828 28444 19717 28472
rect 17828 28432 17834 28444
rect 19705 28441 19717 28444
rect 19751 28441 19763 28475
rect 22940 28472 22968 28571
rect 23216 28540 23244 28639
rect 24688 28617 24716 28648
rect 24762 28636 24768 28648
rect 24820 28676 24826 28688
rect 26160 28676 26188 28704
rect 27632 28676 27660 28716
rect 28077 28713 28089 28747
rect 28123 28744 28135 28747
rect 28166 28744 28172 28756
rect 28123 28716 28172 28744
rect 28123 28713 28135 28716
rect 28077 28707 28135 28713
rect 28166 28704 28172 28716
rect 28224 28704 28230 28756
rect 34057 28747 34115 28753
rect 34057 28713 34069 28747
rect 34103 28744 34115 28747
rect 34790 28744 34796 28756
rect 34103 28716 34796 28744
rect 34103 28713 34115 28716
rect 34057 28707 34115 28713
rect 34790 28704 34796 28716
rect 34848 28704 34854 28756
rect 36725 28747 36783 28753
rect 36725 28713 36737 28747
rect 36771 28744 36783 28747
rect 37366 28744 37372 28756
rect 36771 28716 37372 28744
rect 36771 28713 36783 28716
rect 36725 28707 36783 28713
rect 37366 28704 37372 28716
rect 37424 28704 37430 28756
rect 37458 28704 37464 28756
rect 37516 28744 37522 28756
rect 37737 28747 37795 28753
rect 37737 28744 37749 28747
rect 37516 28716 37749 28744
rect 37516 28704 37522 28716
rect 37737 28713 37749 28716
rect 37783 28713 37795 28747
rect 37737 28707 37795 28713
rect 38381 28747 38439 28753
rect 38381 28713 38393 28747
rect 38427 28744 38439 28747
rect 38562 28744 38568 28756
rect 38427 28716 38568 28744
rect 38427 28713 38439 28716
rect 38381 28707 38439 28713
rect 38562 28704 38568 28716
rect 38620 28704 38626 28756
rect 40126 28704 40132 28756
rect 40184 28744 40190 28756
rect 41049 28747 41107 28753
rect 41049 28744 41061 28747
rect 40184 28716 41061 28744
rect 40184 28704 40190 28716
rect 41049 28713 41061 28716
rect 41095 28713 41107 28747
rect 41049 28707 41107 28713
rect 43993 28747 44051 28753
rect 43993 28713 44005 28747
rect 44039 28744 44051 28747
rect 44082 28744 44088 28756
rect 44039 28716 44088 28744
rect 44039 28713 44051 28716
rect 43993 28707 44051 28713
rect 44082 28704 44088 28716
rect 44140 28744 44146 28756
rect 44542 28744 44548 28756
rect 44140 28716 44548 28744
rect 44140 28704 44146 28716
rect 44542 28704 44548 28716
rect 44600 28704 44606 28756
rect 33686 28676 33692 28688
rect 24820 28648 27568 28676
rect 27632 28648 33692 28676
rect 24820 28636 24826 28648
rect 24673 28611 24731 28617
rect 23860 28580 24532 28608
rect 23860 28549 23888 28580
rect 23661 28543 23719 28549
rect 23661 28540 23673 28543
rect 23216 28512 23673 28540
rect 23661 28509 23673 28512
rect 23707 28509 23719 28543
rect 23661 28503 23719 28509
rect 23845 28543 23903 28549
rect 23845 28509 23857 28543
rect 23891 28509 23903 28543
rect 24397 28543 24455 28549
rect 24397 28540 24409 28543
rect 23845 28503 23903 28509
rect 24320 28512 24409 28540
rect 23750 28472 23756 28484
rect 22940 28444 23756 28472
rect 19705 28435 19763 28441
rect 23750 28432 23756 28444
rect 23808 28432 23814 28484
rect 22094 28404 22100 28416
rect 22055 28376 22100 28404
rect 22094 28364 22100 28376
rect 22152 28364 22158 28416
rect 24320 28404 24348 28512
rect 24397 28509 24409 28512
rect 24443 28509 24455 28543
rect 24504 28540 24532 28580
rect 24673 28577 24685 28611
rect 24719 28577 24731 28611
rect 24673 28571 24731 28577
rect 26142 28568 26148 28620
rect 26200 28608 26206 28620
rect 26421 28611 26479 28617
rect 26421 28608 26433 28611
rect 26200 28580 26433 28608
rect 26200 28568 26206 28580
rect 26421 28577 26433 28580
rect 26467 28577 26479 28611
rect 26421 28571 26479 28577
rect 25314 28540 25320 28552
rect 24504 28512 25320 28540
rect 24397 28503 24455 28509
rect 25314 28500 25320 28512
rect 25372 28540 25378 28552
rect 26050 28540 26056 28552
rect 25372 28512 26056 28540
rect 25372 28500 25378 28512
rect 26050 28500 26056 28512
rect 26108 28500 26114 28552
rect 26326 28540 26332 28552
rect 26287 28512 26332 28540
rect 26326 28500 26332 28512
rect 26384 28500 26390 28552
rect 27430 28540 27436 28552
rect 27391 28512 27436 28540
rect 27430 28500 27436 28512
rect 27488 28500 27494 28552
rect 25961 28475 26019 28481
rect 25961 28441 25973 28475
rect 26007 28472 26019 28475
rect 27448 28472 27476 28500
rect 26007 28444 27476 28472
rect 27540 28472 27568 28648
rect 33686 28636 33692 28648
rect 33744 28636 33750 28688
rect 34698 28636 34704 28688
rect 34756 28676 34762 28688
rect 35253 28679 35311 28685
rect 35253 28676 35265 28679
rect 34756 28648 35265 28676
rect 34756 28636 34762 28648
rect 35253 28645 35265 28648
rect 35299 28645 35311 28679
rect 40494 28676 40500 28688
rect 35253 28639 35311 28645
rect 36832 28648 40500 28676
rect 29454 28608 29460 28620
rect 28368 28580 29460 28608
rect 28368 28549 28396 28580
rect 29454 28568 29460 28580
rect 29512 28568 29518 28620
rect 33502 28568 33508 28620
rect 33560 28608 33566 28620
rect 33965 28611 34023 28617
rect 33965 28608 33977 28611
rect 33560 28580 33977 28608
rect 33560 28568 33566 28580
rect 33965 28577 33977 28580
rect 34011 28577 34023 28611
rect 33965 28571 34023 28577
rect 34149 28611 34207 28617
rect 34149 28577 34161 28611
rect 34195 28608 34207 28611
rect 36832 28608 36860 28648
rect 40494 28636 40500 28648
rect 40552 28636 40558 28688
rect 37826 28608 37832 28620
rect 34195 28580 36860 28608
rect 36924 28580 37832 28608
rect 34195 28577 34207 28580
rect 34149 28571 34207 28577
rect 28353 28543 28411 28549
rect 28353 28509 28365 28543
rect 28399 28509 28411 28543
rect 28353 28503 28411 28509
rect 28445 28543 28503 28549
rect 28445 28509 28457 28543
rect 28491 28509 28503 28543
rect 28445 28503 28503 28509
rect 28460 28472 28488 28503
rect 28534 28500 28540 28552
rect 28592 28540 28598 28552
rect 28592 28512 28637 28540
rect 28592 28500 28598 28512
rect 28718 28500 28724 28552
rect 28776 28540 28782 28552
rect 33870 28540 33876 28552
rect 28776 28512 28821 28540
rect 33831 28512 33876 28540
rect 28776 28500 28782 28512
rect 33870 28500 33876 28512
rect 33928 28500 33934 28552
rect 34701 28543 34759 28549
rect 34701 28540 34713 28543
rect 34164 28512 34713 28540
rect 34164 28484 34192 28512
rect 34701 28509 34713 28512
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 35069 28543 35127 28549
rect 35069 28509 35081 28543
rect 35115 28540 35127 28543
rect 35894 28540 35900 28552
rect 35115 28512 35900 28540
rect 35115 28509 35127 28512
rect 35069 28503 35127 28509
rect 35894 28500 35900 28512
rect 35952 28540 35958 28552
rect 36354 28540 36360 28552
rect 35952 28512 36360 28540
rect 35952 28500 35958 28512
rect 36354 28500 36360 28512
rect 36412 28500 36418 28552
rect 36924 28549 36952 28580
rect 37826 28568 37832 28580
rect 37884 28568 37890 28620
rect 43165 28611 43223 28617
rect 43165 28577 43177 28611
rect 43211 28608 43223 28611
rect 44726 28608 44732 28620
rect 43211 28580 44732 28608
rect 43211 28577 43223 28580
rect 43165 28571 43223 28577
rect 44726 28568 44732 28580
rect 44784 28568 44790 28620
rect 46293 28611 46351 28617
rect 46293 28577 46305 28611
rect 46339 28608 46351 28611
rect 47670 28608 47676 28620
rect 46339 28580 47676 28608
rect 46339 28577 46351 28580
rect 46293 28571 46351 28577
rect 47670 28568 47676 28580
rect 47728 28568 47734 28620
rect 36909 28543 36967 28549
rect 36909 28509 36921 28543
rect 36955 28509 36967 28543
rect 36909 28503 36967 28509
rect 36998 28500 37004 28552
rect 37056 28540 37062 28552
rect 37185 28543 37243 28549
rect 37185 28540 37197 28543
rect 37056 28512 37197 28540
rect 37056 28500 37062 28512
rect 37185 28509 37197 28512
rect 37231 28509 37243 28543
rect 37642 28540 37648 28552
rect 37603 28512 37648 28540
rect 37185 28503 37243 28509
rect 37642 28500 37648 28512
rect 37700 28500 37706 28552
rect 38102 28500 38108 28552
rect 38160 28540 38166 28552
rect 38289 28543 38347 28549
rect 38289 28540 38301 28543
rect 38160 28512 38301 28540
rect 38160 28500 38166 28512
rect 38289 28509 38301 28512
rect 38335 28509 38347 28543
rect 38289 28503 38347 28509
rect 40034 28500 40040 28552
rect 40092 28540 40098 28552
rect 40497 28543 40555 28549
rect 40497 28540 40509 28543
rect 40092 28512 40509 28540
rect 40092 28500 40098 28512
rect 40497 28509 40509 28512
rect 40543 28540 40555 28543
rect 40678 28540 40684 28552
rect 40543 28512 40684 28540
rect 40543 28509 40555 28512
rect 40497 28503 40555 28509
rect 40678 28500 40684 28512
rect 40736 28500 40742 28552
rect 40862 28500 40868 28552
rect 40920 28540 40926 28552
rect 40957 28543 41015 28549
rect 40957 28540 40969 28543
rect 40920 28512 40969 28540
rect 40920 28500 40926 28512
rect 40957 28509 40969 28512
rect 41003 28509 41015 28543
rect 43346 28540 43352 28552
rect 43307 28512 43352 28540
rect 40957 28503 41015 28509
rect 43346 28500 43352 28512
rect 43404 28500 43410 28552
rect 43533 28543 43591 28549
rect 43533 28509 43545 28543
rect 43579 28540 43591 28543
rect 44177 28543 44235 28549
rect 44177 28540 44189 28543
rect 43579 28512 44189 28540
rect 43579 28509 43591 28512
rect 43533 28503 43591 28509
rect 44177 28509 44189 28512
rect 44223 28509 44235 28543
rect 44177 28503 44235 28509
rect 33134 28472 33140 28484
rect 27540 28444 33140 28472
rect 26007 28441 26019 28444
rect 25961 28435 26019 28441
rect 33134 28432 33140 28444
rect 33192 28432 33198 28484
rect 34146 28432 34152 28484
rect 34204 28432 34210 28484
rect 34238 28432 34244 28484
rect 34296 28472 34302 28484
rect 34885 28475 34943 28481
rect 34885 28472 34897 28475
rect 34296 28444 34897 28472
rect 34296 28432 34302 28444
rect 34885 28441 34897 28444
rect 34931 28441 34943 28475
rect 34885 28435 34943 28441
rect 34977 28475 35035 28481
rect 34977 28441 34989 28475
rect 35023 28472 35035 28475
rect 35986 28472 35992 28484
rect 35023 28444 35992 28472
rect 35023 28441 35035 28444
rect 34977 28435 35035 28441
rect 35986 28432 35992 28444
rect 36044 28432 36050 28484
rect 36170 28432 36176 28484
rect 36228 28472 36234 28484
rect 37093 28475 37151 28481
rect 37093 28472 37105 28475
rect 36228 28444 37105 28472
rect 36228 28432 36234 28444
rect 37093 28441 37105 28444
rect 37139 28441 37151 28475
rect 37093 28435 37151 28441
rect 40313 28475 40371 28481
rect 40313 28441 40325 28475
rect 40359 28472 40371 28475
rect 42978 28472 42984 28484
rect 40359 28444 42984 28472
rect 40359 28441 40371 28444
rect 40313 28435 40371 28441
rect 42978 28432 42984 28444
rect 43036 28432 43042 28484
rect 46477 28475 46535 28481
rect 46477 28441 46489 28475
rect 46523 28472 46535 28475
rect 46934 28472 46940 28484
rect 46523 28444 46940 28472
rect 46523 28441 46535 28444
rect 46477 28435 46535 28441
rect 46934 28432 46940 28444
rect 46992 28432 46998 28484
rect 48130 28472 48136 28484
rect 48091 28444 48136 28472
rect 48130 28432 48136 28444
rect 48188 28432 48194 28484
rect 27525 28407 27583 28413
rect 27525 28404 27537 28407
rect 24320 28376 27537 28404
rect 27525 28373 27537 28376
rect 27571 28404 27583 28407
rect 27614 28404 27620 28416
rect 27571 28376 27620 28404
rect 27571 28373 27583 28376
rect 27525 28367 27583 28373
rect 27614 28364 27620 28376
rect 27672 28364 27678 28416
rect 29546 28364 29552 28416
rect 29604 28404 29610 28416
rect 34606 28404 34612 28416
rect 29604 28376 34612 28404
rect 29604 28364 29610 28376
rect 34606 28364 34612 28376
rect 34664 28364 34670 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 16758 28160 16764 28212
rect 16816 28200 16822 28212
rect 17126 28200 17132 28212
rect 16816 28172 17132 28200
rect 16816 28160 16822 28172
rect 17126 28160 17132 28172
rect 17184 28200 17190 28212
rect 22830 28200 22836 28212
rect 17184 28172 18552 28200
rect 22743 28172 22836 28200
rect 17184 28160 17190 28172
rect 18138 28132 18144 28144
rect 18099 28104 18144 28132
rect 18138 28092 18144 28104
rect 18196 28132 18202 28144
rect 18414 28132 18420 28144
rect 18196 28104 18420 28132
rect 18196 28092 18202 28104
rect 18414 28092 18420 28104
rect 18472 28092 18478 28144
rect 18524 28132 18552 28172
rect 22830 28160 22836 28172
rect 22888 28200 22894 28212
rect 23661 28203 23719 28209
rect 23661 28200 23673 28203
rect 22888 28172 23673 28200
rect 22888 28160 22894 28172
rect 23661 28169 23673 28172
rect 23707 28169 23719 28203
rect 23661 28163 23719 28169
rect 26326 28160 26332 28212
rect 26384 28200 26390 28212
rect 27341 28203 27399 28209
rect 27341 28200 27353 28203
rect 26384 28172 27353 28200
rect 26384 28160 26390 28172
rect 27341 28169 27353 28172
rect 27387 28169 27399 28203
rect 27341 28163 27399 28169
rect 27430 28160 27436 28212
rect 27488 28200 27494 28212
rect 28261 28203 28319 28209
rect 28261 28200 28273 28203
rect 27488 28172 28273 28200
rect 27488 28160 27494 28172
rect 28261 28169 28273 28172
rect 28307 28169 28319 28203
rect 28261 28163 28319 28169
rect 28534 28160 28540 28212
rect 28592 28200 28598 28212
rect 28905 28203 28963 28209
rect 28905 28200 28917 28203
rect 28592 28172 28917 28200
rect 28592 28160 28598 28172
rect 28905 28169 28917 28172
rect 28951 28169 28963 28203
rect 28905 28163 28963 28169
rect 31754 28160 31760 28212
rect 31812 28200 31818 28212
rect 32398 28200 32404 28212
rect 31812 28172 32404 28200
rect 31812 28160 31818 28172
rect 32398 28160 32404 28172
rect 32456 28160 32462 28212
rect 33965 28203 34023 28209
rect 33965 28169 33977 28203
rect 34011 28200 34023 28203
rect 34422 28200 34428 28212
rect 34011 28172 34428 28200
rect 34011 28169 34023 28172
rect 33965 28163 34023 28169
rect 34422 28160 34428 28172
rect 34480 28160 34486 28212
rect 35253 28203 35311 28209
rect 35253 28169 35265 28203
rect 35299 28200 35311 28203
rect 35894 28200 35900 28212
rect 35299 28172 35900 28200
rect 35299 28169 35311 28172
rect 35253 28163 35311 28169
rect 35894 28160 35900 28172
rect 35952 28160 35958 28212
rect 40586 28200 40592 28212
rect 40547 28172 40592 28200
rect 40586 28160 40592 28172
rect 40644 28200 40650 28212
rect 41230 28200 41236 28212
rect 40644 28172 41236 28200
rect 40644 28160 40650 28172
rect 41230 28160 41236 28172
rect 41288 28160 41294 28212
rect 45833 28203 45891 28209
rect 45833 28169 45845 28203
rect 45879 28200 45891 28203
rect 46474 28200 46480 28212
rect 45879 28172 46480 28200
rect 45879 28169 45891 28172
rect 45833 28163 45891 28169
rect 46474 28160 46480 28172
rect 46532 28160 46538 28212
rect 31938 28132 31944 28144
rect 18524 28104 31944 28132
rect 31938 28092 31944 28104
rect 31996 28092 32002 28144
rect 32306 28092 32312 28144
rect 32364 28132 32370 28144
rect 43432 28135 43490 28141
rect 32364 28104 32409 28132
rect 40788 28104 41368 28132
rect 32364 28092 32370 28104
rect 40788 28076 40816 28104
rect 17034 28064 17040 28076
rect 16995 28036 17040 28064
rect 17034 28024 17040 28036
rect 17092 28024 17098 28076
rect 17221 28067 17279 28073
rect 17221 28033 17233 28067
rect 17267 28064 17279 28067
rect 17770 28064 17776 28076
rect 17267 28036 17776 28064
rect 17267 28033 17279 28036
rect 17221 28027 17279 28033
rect 17770 28024 17776 28036
rect 17828 28024 17834 28076
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22465 28067 22523 28073
rect 22465 28064 22477 28067
rect 22152 28036 22477 28064
rect 22152 28024 22158 28036
rect 22465 28033 22477 28036
rect 22511 28033 22523 28067
rect 23474 28064 23480 28076
rect 23435 28036 23480 28064
rect 22465 28027 22523 28033
rect 23474 28024 23480 28036
rect 23532 28024 23538 28076
rect 23750 28064 23756 28076
rect 23711 28036 23756 28064
rect 23750 28024 23756 28036
rect 23808 28024 23814 28076
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28064 25651 28067
rect 26142 28064 26148 28076
rect 25639 28036 26148 28064
rect 25639 28033 25651 28036
rect 25593 28027 25651 28033
rect 26142 28024 26148 28036
rect 26200 28024 26206 28076
rect 26418 28024 26424 28076
rect 26476 28064 26482 28076
rect 26973 28067 27031 28073
rect 26973 28064 26985 28067
rect 26476 28036 26985 28064
rect 26476 28024 26482 28036
rect 26973 28033 26985 28036
rect 27019 28033 27031 28067
rect 27154 28064 27160 28076
rect 27115 28036 27160 28064
rect 26973 28027 27031 28033
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 28629 28067 28687 28073
rect 28629 28033 28641 28067
rect 28675 28064 28687 28067
rect 29362 28064 29368 28076
rect 28675 28036 29368 28064
rect 28675 28033 28687 28036
rect 28629 28027 28687 28033
rect 29362 28024 29368 28036
rect 29420 28024 29426 28076
rect 29457 28067 29515 28073
rect 29457 28033 29469 28067
rect 29503 28064 29515 28067
rect 30374 28064 30380 28076
rect 29503 28036 30380 28064
rect 29503 28033 29515 28036
rect 29457 28027 29515 28033
rect 30374 28024 30380 28036
rect 30432 28024 30438 28076
rect 31297 28067 31355 28073
rect 31297 28033 31309 28067
rect 31343 28033 31355 28067
rect 31297 28027 31355 28033
rect 22554 27996 22560 28008
rect 22515 27968 22560 27996
rect 22554 27956 22560 27968
rect 22612 27956 22618 28008
rect 25958 27996 25964 28008
rect 25919 27968 25964 27996
rect 25958 27956 25964 27968
rect 26016 27956 26022 28008
rect 26053 27999 26111 28005
rect 26053 27965 26065 27999
rect 26099 27965 26111 27999
rect 28718 27996 28724 28008
rect 28679 27968 28724 27996
rect 26053 27959 26111 27965
rect 25222 27888 25228 27940
rect 25280 27928 25286 27940
rect 26068 27928 26096 27959
rect 28718 27956 28724 27968
rect 28776 27956 28782 28008
rect 27982 27928 27988 27940
rect 25280 27900 27988 27928
rect 25280 27888 25286 27900
rect 27982 27888 27988 27900
rect 28040 27928 28046 27940
rect 29914 27928 29920 27940
rect 28040 27900 29920 27928
rect 28040 27888 28046 27900
rect 29914 27888 29920 27900
rect 29972 27888 29978 27940
rect 31312 27928 31340 28027
rect 31478 28024 31484 28076
rect 31536 28064 31542 28076
rect 31573 28067 31631 28073
rect 31573 28064 31585 28067
rect 31536 28036 31585 28064
rect 31536 28024 31542 28036
rect 31573 28033 31585 28036
rect 31619 28064 31631 28067
rect 31846 28064 31852 28076
rect 31619 28036 31852 28064
rect 31619 28033 31631 28036
rect 31573 28027 31631 28033
rect 31846 28024 31852 28036
rect 31904 28024 31910 28076
rect 32125 28067 32183 28073
rect 32125 28033 32137 28067
rect 32171 28033 32183 28067
rect 32125 28027 32183 28033
rect 32140 27996 32168 28027
rect 32398 28024 32404 28076
rect 32456 28064 32462 28076
rect 33870 28064 33876 28076
rect 32456 28036 32501 28064
rect 33831 28036 33876 28064
rect 32456 28024 32462 28036
rect 33870 28024 33876 28036
rect 33928 28024 33934 28076
rect 34698 28024 34704 28076
rect 34756 28064 34762 28076
rect 35161 28067 35219 28073
rect 35161 28064 35173 28067
rect 34756 28036 35173 28064
rect 34756 28024 34762 28036
rect 35161 28033 35173 28036
rect 35207 28033 35219 28067
rect 35161 28027 35219 28033
rect 40218 28024 40224 28076
rect 40276 28064 40282 28076
rect 40405 28067 40463 28073
rect 40405 28064 40417 28067
rect 40276 28036 40417 28064
rect 40276 28024 40282 28036
rect 40405 28033 40417 28036
rect 40451 28033 40463 28067
rect 40405 28027 40463 28033
rect 40681 28067 40739 28073
rect 40681 28033 40693 28067
rect 40727 28064 40739 28067
rect 40770 28064 40776 28076
rect 40727 28036 40776 28064
rect 40727 28033 40739 28036
rect 40681 28027 40739 28033
rect 40770 28024 40776 28036
rect 40828 28024 40834 28076
rect 41138 28064 41144 28076
rect 41099 28036 41144 28064
rect 41138 28024 41144 28036
rect 41196 28024 41202 28076
rect 41340 28073 41368 28104
rect 43432 28101 43444 28135
rect 43478 28132 43490 28135
rect 44266 28132 44272 28144
rect 43478 28104 44272 28132
rect 43478 28101 43490 28104
rect 43432 28095 43490 28101
rect 44266 28092 44272 28104
rect 44324 28092 44330 28144
rect 41325 28067 41383 28073
rect 41325 28033 41337 28067
rect 41371 28033 41383 28067
rect 45741 28067 45799 28073
rect 41325 28027 41383 28033
rect 43088 28036 44220 28064
rect 32140 27968 32260 27996
rect 32125 27931 32183 27937
rect 32125 27928 32137 27931
rect 31312 27900 32137 27928
rect 32125 27897 32137 27900
rect 32171 27897 32183 27931
rect 32232 27928 32260 27968
rect 36630 27956 36636 28008
rect 36688 27996 36694 28008
rect 42426 27996 42432 28008
rect 36688 27968 42432 27996
rect 36688 27956 36694 27968
rect 42426 27956 42432 27968
rect 42484 27996 42490 28008
rect 42610 27996 42616 28008
rect 42484 27968 42616 27996
rect 42484 27956 42490 27968
rect 42610 27956 42616 27968
rect 42668 27956 42674 28008
rect 33318 27928 33324 27940
rect 32232 27900 33324 27928
rect 32125 27891 32183 27897
rect 33318 27888 33324 27900
rect 33376 27888 33382 27940
rect 33686 27888 33692 27940
rect 33744 27928 33750 27940
rect 43088 27928 43116 28036
rect 43165 27999 43223 28005
rect 43165 27965 43177 27999
rect 43211 27965 43223 27999
rect 44192 27996 44220 28036
rect 45741 28033 45753 28067
rect 45787 28064 45799 28067
rect 45830 28064 45836 28076
rect 45787 28036 45836 28064
rect 45787 28033 45799 28036
rect 45741 28027 45799 28033
rect 45830 28024 45836 28036
rect 45888 28024 45894 28076
rect 46382 28064 46388 28076
rect 46343 28036 46388 28064
rect 46382 28024 46388 28036
rect 46440 28024 46446 28076
rect 46400 27996 46428 28024
rect 44192 27968 46428 27996
rect 43165 27959 43223 27965
rect 33744 27900 43116 27928
rect 33744 27888 33750 27900
rect 22646 27820 22652 27872
rect 22704 27860 22710 27872
rect 23293 27863 23351 27869
rect 23293 27860 23305 27863
rect 22704 27832 23305 27860
rect 22704 27820 22710 27832
rect 23293 27829 23305 27832
rect 23339 27829 23351 27863
rect 23293 27823 23351 27829
rect 24946 27820 24952 27872
rect 25004 27860 25010 27872
rect 26237 27863 26295 27869
rect 26237 27860 26249 27863
rect 25004 27832 26249 27860
rect 25004 27820 25010 27832
rect 26237 27829 26249 27832
rect 26283 27829 26295 27863
rect 29546 27860 29552 27872
rect 29507 27832 29552 27860
rect 26237 27823 26295 27829
rect 29546 27820 29552 27832
rect 29604 27820 29610 27872
rect 31110 27860 31116 27872
rect 31071 27832 31116 27860
rect 31110 27820 31116 27832
rect 31168 27820 31174 27872
rect 31481 27863 31539 27869
rect 31481 27829 31493 27863
rect 31527 27860 31539 27863
rect 33134 27860 33140 27872
rect 31527 27832 33140 27860
rect 31527 27829 31539 27832
rect 31481 27823 31539 27829
rect 33134 27820 33140 27832
rect 33192 27820 33198 27872
rect 40405 27863 40463 27869
rect 40405 27829 40417 27863
rect 40451 27860 40463 27863
rect 40586 27860 40592 27872
rect 40451 27832 40592 27860
rect 40451 27829 40463 27832
rect 40405 27823 40463 27829
rect 40586 27820 40592 27832
rect 40644 27820 40650 27872
rect 41141 27863 41199 27869
rect 41141 27829 41153 27863
rect 41187 27860 41199 27863
rect 41506 27860 41512 27872
rect 41187 27832 41512 27860
rect 41187 27829 41199 27832
rect 41141 27823 41199 27829
rect 41506 27820 41512 27832
rect 41564 27820 41570 27872
rect 43180 27860 43208 27959
rect 43806 27860 43812 27872
rect 43180 27832 43812 27860
rect 43806 27820 43812 27832
rect 43864 27820 43870 27872
rect 44545 27863 44603 27869
rect 44545 27829 44557 27863
rect 44591 27860 44603 27863
rect 45278 27860 45284 27872
rect 44591 27832 45284 27860
rect 44591 27829 44603 27832
rect 44545 27823 44603 27829
rect 45278 27820 45284 27832
rect 45336 27820 45342 27872
rect 46474 27860 46480 27872
rect 46435 27832 46480 27860
rect 46474 27820 46480 27832
rect 46532 27820 46538 27872
rect 47762 27860 47768 27872
rect 47723 27832 47768 27860
rect 47762 27820 47768 27832
rect 47820 27820 47826 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 26142 27656 26148 27668
rect 26103 27628 26148 27656
rect 26142 27616 26148 27628
rect 26200 27616 26206 27668
rect 28718 27616 28724 27668
rect 28776 27656 28782 27668
rect 28905 27659 28963 27665
rect 28905 27656 28917 27659
rect 28776 27628 28917 27656
rect 28776 27616 28782 27628
rect 28905 27625 28917 27628
rect 28951 27625 28963 27659
rect 28905 27619 28963 27625
rect 33965 27659 34023 27665
rect 33965 27625 33977 27659
rect 34011 27656 34023 27659
rect 34238 27656 34244 27668
rect 34011 27628 34244 27656
rect 34011 27625 34023 27628
rect 33965 27619 34023 27625
rect 34238 27616 34244 27628
rect 34296 27616 34302 27668
rect 37642 27616 37648 27668
rect 37700 27656 37706 27668
rect 38289 27659 38347 27665
rect 38289 27656 38301 27659
rect 37700 27628 38301 27656
rect 37700 27616 37706 27628
rect 38289 27625 38301 27628
rect 38335 27625 38347 27659
rect 40037 27659 40095 27665
rect 38289 27619 38347 27625
rect 38396 27628 39160 27656
rect 23750 27548 23756 27600
rect 23808 27588 23814 27600
rect 24949 27591 25007 27597
rect 24949 27588 24961 27591
rect 23808 27560 24961 27588
rect 23808 27548 23814 27560
rect 24949 27557 24961 27560
rect 24995 27557 25007 27591
rect 26050 27588 26056 27600
rect 24949 27551 25007 27557
rect 25240 27560 26056 27588
rect 25240 27529 25268 27560
rect 26050 27548 26056 27560
rect 26108 27588 26114 27600
rect 26418 27588 26424 27600
rect 26108 27560 26424 27588
rect 26108 27548 26114 27560
rect 26418 27548 26424 27560
rect 26476 27548 26482 27600
rect 26510 27548 26516 27600
rect 26568 27588 26574 27600
rect 26568 27560 29316 27588
rect 26568 27548 26574 27560
rect 25225 27523 25283 27529
rect 25225 27489 25237 27523
rect 25271 27489 25283 27523
rect 25225 27483 25283 27489
rect 25317 27523 25375 27529
rect 25317 27489 25329 27523
rect 25363 27520 25375 27523
rect 25498 27520 25504 27532
rect 25363 27492 25504 27520
rect 25363 27489 25375 27492
rect 25317 27483 25375 27489
rect 25498 27480 25504 27492
rect 25556 27480 25562 27532
rect 29288 27520 29316 27560
rect 29362 27548 29368 27600
rect 29420 27588 29426 27600
rect 29917 27591 29975 27597
rect 29917 27588 29929 27591
rect 29420 27560 29929 27588
rect 29420 27548 29426 27560
rect 29917 27557 29929 27560
rect 29963 27557 29975 27591
rect 29917 27551 29975 27557
rect 34606 27548 34612 27600
rect 34664 27588 34670 27600
rect 38396 27588 38424 27628
rect 34664 27560 38424 27588
rect 38473 27591 38531 27597
rect 34664 27548 34670 27560
rect 29288 27492 29868 27520
rect 8386 27412 8392 27464
rect 8444 27452 8450 27464
rect 15933 27455 15991 27461
rect 15933 27452 15945 27455
rect 8444 27424 15945 27452
rect 8444 27412 8450 27424
rect 15933 27421 15945 27424
rect 15979 27452 15991 27455
rect 17034 27452 17040 27464
rect 15979 27424 17040 27452
rect 15979 27421 15991 27424
rect 15933 27415 15991 27421
rect 17034 27412 17040 27424
rect 17092 27412 17098 27464
rect 18046 27452 18052 27464
rect 17144 27424 18052 27452
rect 16117 27387 16175 27393
rect 16117 27353 16129 27387
rect 16163 27384 16175 27387
rect 16577 27387 16635 27393
rect 16577 27384 16589 27387
rect 16163 27356 16589 27384
rect 16163 27353 16175 27356
rect 16117 27347 16175 27353
rect 16577 27353 16589 27356
rect 16623 27384 16635 27387
rect 17144 27384 17172 27424
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 25130 27452 25136 27464
rect 25091 27424 25136 27452
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27452 25467 27455
rect 25590 27452 25596 27464
rect 25455 27424 25596 27452
rect 25455 27421 25467 27424
rect 25409 27415 25467 27421
rect 25590 27412 25596 27424
rect 25648 27412 25654 27464
rect 26050 27412 26056 27464
rect 26108 27452 26114 27464
rect 26237 27455 26295 27461
rect 26108 27424 26153 27452
rect 26108 27412 26114 27424
rect 26237 27421 26249 27455
rect 26283 27452 26295 27455
rect 27154 27452 27160 27464
rect 26283 27424 27160 27452
rect 26283 27421 26295 27424
rect 26237 27415 26295 27421
rect 17310 27384 17316 27396
rect 16623 27356 17172 27384
rect 17271 27356 17316 27384
rect 16623 27353 16635 27356
rect 16577 27347 16635 27353
rect 17310 27344 17316 27356
rect 17368 27344 17374 27396
rect 18598 27384 18604 27396
rect 18511 27356 18604 27384
rect 18598 27344 18604 27356
rect 18656 27384 18662 27396
rect 24118 27384 24124 27396
rect 18656 27356 24124 27384
rect 18656 27344 18662 27356
rect 24118 27344 24124 27356
rect 24176 27344 24182 27396
rect 25498 27276 25504 27328
rect 25556 27316 25562 27328
rect 26252 27316 26280 27415
rect 27154 27412 27160 27424
rect 27212 27412 27218 27464
rect 28813 27455 28871 27461
rect 28813 27421 28825 27455
rect 28859 27421 28871 27455
rect 28813 27415 28871 27421
rect 28626 27344 28632 27396
rect 28684 27384 28690 27396
rect 28828 27384 28856 27415
rect 28902 27412 28908 27464
rect 28960 27452 28966 27464
rect 28997 27455 29055 27461
rect 28997 27452 29009 27455
rect 28960 27424 29009 27452
rect 28960 27412 28966 27424
rect 28997 27421 29009 27424
rect 29043 27421 29055 27455
rect 28997 27415 29055 27421
rect 29549 27387 29607 27393
rect 29549 27384 29561 27387
rect 28684 27356 29561 27384
rect 28684 27344 28690 27356
rect 29549 27353 29561 27356
rect 29595 27353 29607 27387
rect 29549 27347 29607 27353
rect 29733 27387 29791 27393
rect 29733 27353 29745 27387
rect 29779 27353 29791 27387
rect 29733 27347 29791 27353
rect 25556 27288 26280 27316
rect 25556 27276 25562 27288
rect 28902 27276 28908 27328
rect 28960 27316 28966 27328
rect 29748 27316 29776 27347
rect 28960 27288 29776 27316
rect 29840 27316 29868 27492
rect 34422 27480 34428 27532
rect 34480 27520 34486 27532
rect 34992 27529 35020 27560
rect 38473 27557 38485 27591
rect 38519 27557 38531 27591
rect 38473 27551 38531 27557
rect 34793 27523 34851 27529
rect 34793 27520 34805 27523
rect 34480 27492 34805 27520
rect 34480 27480 34486 27492
rect 34793 27489 34805 27492
rect 34839 27489 34851 27523
rect 34793 27483 34851 27489
rect 34977 27523 35035 27529
rect 34977 27489 34989 27523
rect 35023 27489 35035 27523
rect 37366 27520 37372 27532
rect 34977 27483 35035 27489
rect 35636 27492 37372 27520
rect 35636 27464 35664 27492
rect 37366 27480 37372 27492
rect 37424 27480 37430 27532
rect 37461 27523 37519 27529
rect 37461 27489 37473 27523
rect 37507 27520 37519 27523
rect 37642 27520 37648 27532
rect 37507 27492 37648 27520
rect 37507 27489 37519 27492
rect 37461 27483 37519 27489
rect 37642 27480 37648 27492
rect 37700 27480 37706 27532
rect 30837 27455 30895 27461
rect 30837 27421 30849 27455
rect 30883 27452 30895 27455
rect 32950 27452 32956 27464
rect 30883 27424 32956 27452
rect 30883 27421 30895 27424
rect 30837 27415 30895 27421
rect 32950 27412 32956 27424
rect 33008 27412 33014 27464
rect 33686 27412 33692 27464
rect 33744 27452 33750 27464
rect 33873 27455 33931 27461
rect 33873 27452 33885 27455
rect 33744 27424 33885 27452
rect 33744 27412 33750 27424
rect 33873 27421 33885 27424
rect 33919 27421 33931 27455
rect 34698 27452 34704 27464
rect 34659 27424 34704 27452
rect 33873 27415 33931 27421
rect 34698 27412 34704 27424
rect 34756 27412 34762 27464
rect 35437 27455 35495 27461
rect 35437 27452 35449 27455
rect 34992 27424 35449 27452
rect 31110 27393 31116 27396
rect 31104 27384 31116 27393
rect 31071 27356 31116 27384
rect 31104 27347 31116 27356
rect 31110 27344 31116 27347
rect 31168 27344 31174 27396
rect 34882 27384 34888 27396
rect 31726 27356 34888 27384
rect 31726 27316 31754 27356
rect 34882 27344 34888 27356
rect 34940 27344 34946 27396
rect 34992 27393 35020 27424
rect 35437 27421 35449 27424
rect 35483 27421 35495 27455
rect 35618 27452 35624 27464
rect 35579 27424 35624 27452
rect 35437 27415 35495 27421
rect 35618 27412 35624 27424
rect 35676 27412 35682 27464
rect 37185 27455 37243 27461
rect 37185 27421 37197 27455
rect 37231 27452 37243 27455
rect 37274 27452 37280 27464
rect 37231 27424 37280 27452
rect 37231 27421 37243 27424
rect 37185 27415 37243 27421
rect 37274 27412 37280 27424
rect 37332 27412 37338 27464
rect 38488 27452 38516 27551
rect 38562 27548 38568 27600
rect 38620 27588 38626 27600
rect 38620 27560 39068 27588
rect 38620 27548 38626 27560
rect 39040 27529 39068 27560
rect 39025 27523 39083 27529
rect 39025 27489 39037 27523
rect 39071 27489 39083 27523
rect 39132 27520 39160 27628
rect 40037 27625 40049 27659
rect 40083 27656 40095 27659
rect 41138 27656 41144 27668
rect 40083 27628 41144 27656
rect 40083 27625 40095 27628
rect 40037 27619 40095 27625
rect 41138 27616 41144 27628
rect 41196 27616 41202 27668
rect 39482 27548 39488 27600
rect 39540 27588 39546 27600
rect 39945 27591 40003 27597
rect 39945 27588 39957 27591
rect 39540 27560 39957 27588
rect 39540 27548 39546 27560
rect 39945 27557 39957 27560
rect 39991 27588 40003 27591
rect 47762 27588 47768 27600
rect 39991 27560 40816 27588
rect 39991 27557 40003 27560
rect 39945 27551 40003 27557
rect 39206 27520 39212 27532
rect 39132 27492 39212 27520
rect 39025 27483 39083 27489
rect 39206 27480 39212 27492
rect 39264 27480 39270 27532
rect 39390 27480 39396 27532
rect 39448 27520 39454 27532
rect 40129 27523 40187 27529
rect 40129 27520 40141 27523
rect 39448 27492 40141 27520
rect 39448 27480 39454 27492
rect 40129 27489 40141 27492
rect 40175 27489 40187 27523
rect 40129 27483 40187 27489
rect 38933 27455 38991 27461
rect 38933 27452 38945 27455
rect 37384 27424 38240 27452
rect 38488 27424 38945 27452
rect 34977 27387 35035 27393
rect 34977 27353 34989 27387
rect 35023 27353 35035 27387
rect 37384 27384 37412 27424
rect 38102 27384 38108 27396
rect 34977 27347 35035 27353
rect 35360 27356 37412 27384
rect 38063 27356 38108 27384
rect 29840 27288 31754 27316
rect 28960 27276 28966 27288
rect 31846 27276 31852 27328
rect 31904 27316 31910 27328
rect 32214 27316 32220 27328
rect 31904 27288 32220 27316
rect 31904 27276 31910 27288
rect 32214 27276 32220 27288
rect 32272 27276 32278 27328
rect 33134 27276 33140 27328
rect 33192 27316 33198 27328
rect 35360 27316 35388 27356
rect 38102 27344 38108 27356
rect 38160 27344 38166 27396
rect 38212 27384 38240 27424
rect 38933 27421 38945 27424
rect 38979 27452 38991 27455
rect 39482 27452 39488 27464
rect 38979 27424 39488 27452
rect 38979 27421 38991 27424
rect 38933 27415 38991 27421
rect 39482 27412 39488 27424
rect 39540 27412 39546 27464
rect 40788 27461 40816 27560
rect 46308 27560 47768 27588
rect 46308 27529 46336 27560
rect 47762 27548 47768 27560
rect 47820 27548 47826 27600
rect 46293 27523 46351 27529
rect 46293 27489 46305 27523
rect 46339 27489 46351 27523
rect 46474 27520 46480 27532
rect 46435 27492 46480 27520
rect 46293 27483 46351 27489
rect 46474 27480 46480 27492
rect 46532 27480 46538 27532
rect 46842 27520 46848 27532
rect 46803 27492 46848 27520
rect 46842 27480 46848 27492
rect 46900 27480 46906 27532
rect 39853 27455 39911 27461
rect 39853 27421 39865 27455
rect 39899 27452 39911 27455
rect 40681 27455 40739 27461
rect 40681 27452 40693 27455
rect 39899 27424 40693 27452
rect 39899 27421 39911 27424
rect 39853 27415 39911 27421
rect 40681 27421 40693 27424
rect 40727 27421 40739 27455
rect 40681 27415 40739 27421
rect 40773 27455 40831 27461
rect 40773 27421 40785 27455
rect 40819 27421 40831 27455
rect 40773 27415 40831 27421
rect 41417 27455 41475 27461
rect 41417 27421 41429 27455
rect 41463 27452 41475 27455
rect 43806 27452 43812 27464
rect 41463 27424 43812 27452
rect 41463 27421 41475 27424
rect 41417 27415 41475 27421
rect 39209 27387 39267 27393
rect 39209 27384 39221 27387
rect 38212 27356 39221 27384
rect 39209 27353 39221 27356
rect 39255 27384 39267 27387
rect 40310 27384 40316 27396
rect 39255 27356 40316 27384
rect 39255 27353 39267 27356
rect 39209 27347 39267 27353
rect 40310 27344 40316 27356
rect 40368 27344 40374 27396
rect 40696 27384 40724 27415
rect 43806 27412 43812 27424
rect 43864 27412 43870 27464
rect 40862 27384 40868 27396
rect 40696 27356 40868 27384
rect 40862 27344 40868 27356
rect 40920 27384 40926 27396
rect 40920 27356 41092 27384
rect 40920 27344 40926 27356
rect 35526 27316 35532 27328
rect 33192 27288 35388 27316
rect 35487 27288 35532 27316
rect 33192 27276 33198 27288
rect 35526 27276 35532 27288
rect 35584 27276 35590 27328
rect 36998 27316 37004 27328
rect 36959 27288 37004 27316
rect 36998 27276 37004 27288
rect 37056 27276 37062 27328
rect 37366 27276 37372 27328
rect 37424 27316 37430 27328
rect 38305 27319 38363 27325
rect 38305 27316 38317 27319
rect 37424 27288 38317 27316
rect 37424 27276 37430 27288
rect 38305 27285 38317 27288
rect 38351 27316 38363 27319
rect 38470 27316 38476 27328
rect 38351 27288 38476 27316
rect 38351 27285 38363 27288
rect 38305 27279 38363 27285
rect 38470 27276 38476 27288
rect 38528 27276 38534 27328
rect 38562 27276 38568 27328
rect 38620 27316 38626 27328
rect 38933 27319 38991 27325
rect 38933 27316 38945 27319
rect 38620 27288 38945 27316
rect 38620 27276 38626 27288
rect 38933 27285 38945 27288
rect 38979 27285 38991 27319
rect 38933 27279 38991 27285
rect 40770 27276 40776 27328
rect 40828 27316 40834 27328
rect 40957 27319 41015 27325
rect 40957 27316 40969 27319
rect 40828 27288 40969 27316
rect 40828 27276 40834 27288
rect 40957 27285 40969 27288
rect 41003 27285 41015 27319
rect 41064 27316 41092 27356
rect 41506 27344 41512 27396
rect 41564 27384 41570 27396
rect 41662 27387 41720 27393
rect 41662 27384 41674 27387
rect 41564 27356 41674 27384
rect 41564 27344 41570 27356
rect 41662 27353 41674 27356
rect 41708 27353 41720 27387
rect 41662 27347 41720 27353
rect 42886 27344 42892 27396
rect 42944 27384 42950 27396
rect 43349 27387 43407 27393
rect 43349 27384 43361 27387
rect 42944 27356 43361 27384
rect 42944 27344 42950 27356
rect 43349 27353 43361 27356
rect 43395 27384 43407 27387
rect 46014 27384 46020 27396
rect 43395 27356 46020 27384
rect 43395 27353 43407 27356
rect 43349 27347 43407 27353
rect 46014 27344 46020 27356
rect 46072 27344 46078 27396
rect 42797 27319 42855 27325
rect 42797 27316 42809 27319
rect 41064 27288 42809 27316
rect 40957 27279 41015 27285
rect 42797 27285 42809 27288
rect 42843 27285 42855 27319
rect 43438 27316 43444 27328
rect 43399 27288 43444 27316
rect 42797 27279 42855 27285
rect 43438 27276 43444 27288
rect 43496 27276 43502 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 16942 27072 16948 27124
rect 17000 27072 17006 27124
rect 17034 27072 17040 27124
rect 17092 27112 17098 27124
rect 42889 27115 42947 27121
rect 17092 27084 41414 27112
rect 17092 27072 17098 27084
rect 7837 27047 7895 27053
rect 7837 27013 7849 27047
rect 7883 27044 7895 27047
rect 8386 27044 8392 27056
rect 7883 27016 8392 27044
rect 7883 27013 7895 27016
rect 7837 27007 7895 27013
rect 8386 27004 8392 27016
rect 8444 27004 8450 27056
rect 16960 27044 16988 27072
rect 18325 27047 18383 27053
rect 18325 27044 18337 27047
rect 16960 27016 18337 27044
rect 18325 27013 18337 27016
rect 18371 27044 18383 27047
rect 21910 27044 21916 27056
rect 18371 27016 21916 27044
rect 18371 27013 18383 27016
rect 18325 27007 18383 27013
rect 21910 27004 21916 27016
rect 21968 27004 21974 27056
rect 25406 27004 25412 27056
rect 25464 27044 25470 27056
rect 34416 27047 34474 27053
rect 25464 27016 34284 27044
rect 25464 27004 25470 27016
rect 16666 26936 16672 26988
rect 16724 26976 16730 26988
rect 16945 26979 17003 26985
rect 16945 26976 16957 26979
rect 16724 26948 16957 26976
rect 16724 26936 16730 26948
rect 16945 26945 16957 26948
rect 16991 26976 17003 26979
rect 18046 26976 18052 26988
rect 16991 26948 18052 26976
rect 16991 26945 17003 26948
rect 16945 26939 17003 26945
rect 18046 26936 18052 26948
rect 18104 26936 18110 26988
rect 23201 26979 23259 26985
rect 23201 26945 23213 26979
rect 23247 26945 23259 26979
rect 23201 26939 23259 26945
rect 24765 26979 24823 26985
rect 24765 26945 24777 26979
rect 24811 26976 24823 26979
rect 25130 26976 25136 26988
rect 24811 26948 25136 26976
rect 24811 26945 24823 26948
rect 24765 26939 24823 26945
rect 17497 26911 17555 26917
rect 17497 26877 17509 26911
rect 17543 26908 17555 26911
rect 17862 26908 17868 26920
rect 17543 26880 17868 26908
rect 17543 26877 17555 26880
rect 17497 26871 17555 26877
rect 17862 26868 17868 26880
rect 17920 26868 17926 26920
rect 22554 26868 22560 26920
rect 22612 26908 22618 26920
rect 23014 26908 23020 26920
rect 22612 26880 23020 26908
rect 22612 26868 22618 26880
rect 23014 26868 23020 26880
rect 23072 26908 23078 26920
rect 23109 26911 23167 26917
rect 23109 26908 23121 26911
rect 23072 26880 23121 26908
rect 23072 26868 23078 26880
rect 23109 26877 23121 26880
rect 23155 26877 23167 26911
rect 23109 26871 23167 26877
rect 7926 26772 7932 26784
rect 7887 26744 7932 26772
rect 7926 26732 7932 26744
rect 7984 26732 7990 26784
rect 23216 26772 23244 26939
rect 23569 26843 23627 26849
rect 23569 26809 23581 26843
rect 23615 26840 23627 26843
rect 24780 26840 24808 26939
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 26053 26979 26111 26985
rect 26053 26945 26065 26979
rect 26099 26976 26111 26979
rect 26786 26976 26792 26988
rect 26099 26948 26792 26976
rect 26099 26945 26111 26948
rect 26053 26939 26111 26945
rect 26786 26936 26792 26948
rect 26844 26936 26850 26988
rect 27433 26979 27491 26985
rect 27433 26945 27445 26979
rect 27479 26976 27491 26979
rect 28258 26976 28264 26988
rect 27479 26948 28264 26976
rect 27479 26945 27491 26948
rect 27433 26939 27491 26945
rect 28258 26936 28264 26948
rect 28316 26936 28322 26988
rect 28626 26976 28632 26988
rect 28587 26948 28632 26976
rect 28626 26936 28632 26948
rect 28684 26936 28690 26988
rect 28721 26979 28779 26985
rect 28721 26945 28733 26979
rect 28767 26976 28779 26979
rect 28902 26976 28908 26988
rect 28767 26948 28908 26976
rect 28767 26945 28779 26948
rect 28721 26939 28779 26945
rect 28902 26936 28908 26948
rect 28960 26936 28966 26988
rect 32861 26979 32919 26985
rect 32861 26945 32873 26979
rect 32907 26945 32919 26979
rect 32861 26939 32919 26945
rect 24857 26911 24915 26917
rect 24857 26877 24869 26911
rect 24903 26908 24915 26911
rect 24946 26908 24952 26920
rect 24903 26880 24952 26908
rect 24903 26877 24915 26880
rect 24857 26871 24915 26877
rect 24946 26868 24952 26880
rect 25004 26868 25010 26920
rect 25774 26868 25780 26920
rect 25832 26908 25838 26920
rect 25961 26911 26019 26917
rect 25961 26908 25973 26911
rect 25832 26880 25973 26908
rect 25832 26868 25838 26880
rect 25961 26877 25973 26880
rect 26007 26908 26019 26911
rect 26007 26880 26556 26908
rect 26007 26877 26019 26880
rect 25961 26871 26019 26877
rect 25130 26840 25136 26852
rect 23615 26812 24808 26840
rect 25091 26812 25136 26840
rect 23615 26809 23627 26812
rect 23569 26803 23627 26809
rect 25130 26800 25136 26812
rect 25188 26800 25194 26852
rect 26418 26840 26424 26852
rect 26379 26812 26424 26840
rect 26418 26800 26424 26812
rect 26476 26800 26482 26852
rect 26528 26840 26556 26880
rect 27154 26868 27160 26920
rect 27212 26908 27218 26920
rect 28353 26911 28411 26917
rect 28353 26908 28365 26911
rect 27212 26880 28365 26908
rect 27212 26868 27218 26880
rect 28353 26877 28365 26880
rect 28399 26877 28411 26911
rect 28534 26908 28540 26920
rect 28495 26880 28540 26908
rect 28353 26871 28411 26877
rect 28534 26868 28540 26880
rect 28592 26868 28598 26920
rect 28813 26911 28871 26917
rect 28813 26877 28825 26911
rect 28859 26877 28871 26911
rect 32876 26908 32904 26939
rect 32950 26936 32956 26988
rect 33008 26976 33014 26988
rect 34149 26979 34207 26985
rect 34149 26976 34161 26979
rect 33008 26948 34161 26976
rect 33008 26936 33014 26948
rect 34149 26945 34161 26948
rect 34195 26945 34207 26979
rect 34256 26976 34284 27016
rect 34416 27013 34428 27047
rect 34462 27044 34474 27047
rect 35526 27044 35532 27056
rect 34462 27016 35532 27044
rect 34462 27013 34474 27016
rect 34416 27007 34474 27013
rect 35526 27004 35532 27016
rect 35584 27004 35590 27056
rect 37461 27047 37519 27053
rect 37461 27013 37473 27047
rect 37507 27044 37519 27047
rect 37642 27044 37648 27056
rect 37507 27016 37648 27044
rect 37507 27013 37519 27016
rect 37461 27007 37519 27013
rect 37642 27004 37648 27016
rect 37700 27004 37706 27056
rect 41386 27044 41414 27084
rect 42889 27081 42901 27115
rect 42935 27112 42947 27115
rect 43346 27112 43352 27124
rect 42935 27084 43352 27112
rect 42935 27081 42947 27084
rect 42889 27075 42947 27081
rect 43346 27072 43352 27084
rect 43404 27072 43410 27124
rect 46934 27112 46940 27124
rect 46895 27084 46940 27112
rect 46934 27072 46940 27084
rect 46992 27072 46998 27124
rect 44082 27053 44088 27056
rect 44076 27044 44088 27053
rect 38028 27016 38792 27044
rect 41386 27016 43024 27044
rect 44043 27016 44088 27044
rect 34256 26948 35204 26976
rect 34149 26939 34207 26945
rect 32876 26880 33088 26908
rect 28813 26871 28871 26877
rect 27617 26843 27675 26849
rect 27617 26840 27629 26843
rect 26528 26812 27629 26840
rect 27617 26809 27629 26812
rect 27663 26809 27675 26843
rect 27617 26803 27675 26809
rect 28442 26800 28448 26852
rect 28500 26840 28506 26852
rect 28828 26840 28856 26871
rect 28500 26812 28856 26840
rect 28500 26800 28506 26812
rect 32674 26800 32680 26852
rect 32732 26840 32738 26852
rect 32953 26843 33011 26849
rect 32953 26840 32965 26843
rect 32732 26812 32965 26840
rect 32732 26800 32738 26812
rect 32953 26809 32965 26812
rect 32999 26809 33011 26843
rect 32953 26803 33011 26809
rect 27062 26772 27068 26784
rect 23216 26744 27068 26772
rect 27062 26732 27068 26744
rect 27120 26732 27126 26784
rect 32858 26772 32864 26784
rect 32819 26744 32864 26772
rect 32858 26732 32864 26744
rect 32916 26732 32922 26784
rect 33060 26772 33088 26880
rect 33134 26868 33140 26920
rect 33192 26908 33198 26920
rect 35176 26908 35204 26948
rect 36538 26936 36544 26988
rect 36596 26976 36602 26988
rect 37277 26979 37335 26985
rect 37277 26976 37289 26979
rect 36596 26948 37289 26976
rect 36596 26936 36602 26948
rect 37277 26945 37289 26948
rect 37323 26945 37335 26979
rect 37277 26939 37335 26945
rect 37366 26936 37372 26988
rect 37424 26976 37430 26988
rect 37553 26979 37611 26985
rect 37553 26976 37565 26979
rect 37424 26948 37565 26976
rect 37424 26936 37430 26948
rect 37553 26945 37565 26948
rect 37599 26945 37611 26979
rect 37553 26939 37611 26945
rect 37826 26936 37832 26988
rect 37884 26976 37890 26988
rect 38028 26985 38056 27016
rect 38764 26988 38792 27016
rect 38013 26979 38071 26985
rect 38013 26976 38025 26979
rect 37884 26948 38025 26976
rect 37884 26936 37890 26948
rect 38013 26945 38025 26948
rect 38059 26945 38071 26979
rect 38013 26939 38071 26945
rect 38280 26979 38338 26985
rect 38280 26945 38292 26979
rect 38326 26976 38338 26979
rect 38562 26976 38568 26988
rect 38326 26948 38568 26976
rect 38326 26945 38338 26948
rect 38280 26939 38338 26945
rect 38562 26936 38568 26948
rect 38620 26936 38626 26988
rect 38746 26936 38752 26988
rect 38804 26976 38810 26988
rect 39850 26976 39856 26988
rect 38804 26948 39856 26976
rect 38804 26936 38810 26948
rect 39850 26936 39856 26948
rect 39908 26936 39914 26988
rect 40120 26979 40178 26985
rect 40120 26945 40132 26979
rect 40166 26976 40178 26979
rect 40402 26976 40408 26988
rect 40166 26948 40408 26976
rect 40166 26945 40178 26948
rect 40120 26939 40178 26945
rect 40402 26936 40408 26948
rect 40460 26936 40466 26988
rect 40678 26936 40684 26988
rect 40736 26976 40742 26988
rect 41598 26976 41604 26988
rect 40736 26948 41604 26976
rect 40736 26936 40742 26948
rect 41598 26936 41604 26948
rect 41656 26936 41662 26988
rect 42797 26979 42855 26985
rect 42797 26945 42809 26979
rect 42843 26976 42855 26979
rect 42886 26976 42892 26988
rect 42843 26948 42892 26976
rect 42843 26945 42855 26948
rect 42797 26939 42855 26945
rect 42886 26936 42892 26948
rect 42944 26936 42950 26988
rect 42996 26976 43024 27016
rect 44076 27007 44088 27016
rect 44082 27004 44088 27007
rect 44140 27004 44146 27056
rect 45925 26979 45983 26985
rect 45925 26976 45937 26979
rect 42996 26948 45937 26976
rect 45925 26945 45937 26948
rect 45971 26976 45983 26979
rect 46106 26976 46112 26988
rect 45971 26948 46112 26976
rect 45971 26945 45983 26948
rect 45925 26939 45983 26945
rect 46106 26936 46112 26948
rect 46164 26936 46170 26988
rect 46845 26979 46903 26985
rect 46845 26945 46857 26979
rect 46891 26976 46903 26979
rect 47578 26976 47584 26988
rect 46891 26948 47584 26976
rect 46891 26945 46903 26948
rect 46845 26939 46903 26945
rect 37642 26908 37648 26920
rect 33192 26880 33237 26908
rect 35176 26880 37648 26908
rect 33192 26868 33198 26880
rect 37642 26868 37648 26880
rect 37700 26868 37706 26920
rect 43806 26908 43812 26920
rect 43767 26880 43812 26908
rect 43806 26868 43812 26880
rect 43864 26868 43870 26920
rect 45370 26868 45376 26920
rect 45428 26908 45434 26920
rect 46860 26908 46888 26939
rect 47578 26936 47584 26948
rect 47636 26936 47642 26988
rect 47670 26936 47676 26988
rect 47728 26976 47734 26988
rect 47765 26979 47823 26985
rect 47765 26976 47777 26979
rect 47728 26948 47777 26976
rect 47728 26936 47734 26948
rect 47765 26945 47777 26948
rect 47811 26945 47823 26979
rect 47765 26939 47823 26945
rect 45428 26880 46888 26908
rect 45428 26868 45434 26880
rect 35158 26800 35164 26852
rect 35216 26840 35222 26852
rect 37274 26840 37280 26852
rect 35216 26812 35664 26840
rect 37235 26812 37280 26840
rect 35216 26800 35222 26812
rect 34422 26772 34428 26784
rect 33060 26744 34428 26772
rect 34422 26732 34428 26744
rect 34480 26732 34486 26784
rect 34790 26732 34796 26784
rect 34848 26772 34854 26784
rect 35529 26775 35587 26781
rect 35529 26772 35541 26775
rect 34848 26744 35541 26772
rect 34848 26732 34854 26744
rect 35529 26741 35541 26744
rect 35575 26741 35587 26775
rect 35636 26772 35664 26812
rect 37274 26800 37280 26812
rect 37332 26800 37338 26852
rect 41230 26840 41236 26852
rect 41191 26812 41236 26840
rect 41230 26800 41236 26812
rect 41288 26800 41294 26852
rect 38010 26772 38016 26784
rect 35636 26744 38016 26772
rect 35529 26735 35587 26741
rect 38010 26732 38016 26744
rect 38068 26732 38074 26784
rect 38194 26732 38200 26784
rect 38252 26772 38258 26784
rect 39393 26775 39451 26781
rect 39393 26772 39405 26775
rect 38252 26744 39405 26772
rect 38252 26732 38258 26744
rect 39393 26741 39405 26744
rect 39439 26741 39451 26775
rect 39393 26735 39451 26741
rect 45189 26775 45247 26781
rect 45189 26741 45201 26775
rect 45235 26772 45247 26775
rect 45738 26772 45744 26784
rect 45235 26744 45744 26772
rect 45235 26741 45247 26744
rect 45189 26735 45247 26741
rect 45738 26732 45744 26744
rect 45796 26732 45802 26784
rect 46017 26775 46075 26781
rect 46017 26741 46029 26775
rect 46063 26772 46075 26775
rect 46290 26772 46296 26784
rect 46063 26744 46296 26772
rect 46063 26741 46075 26744
rect 46017 26735 46075 26741
rect 46290 26732 46296 26744
rect 46348 26732 46354 26784
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 8202 26528 8208 26580
rect 8260 26568 8266 26580
rect 25406 26568 25412 26580
rect 8260 26540 25412 26568
rect 8260 26528 8266 26540
rect 25406 26528 25412 26540
rect 25464 26528 25470 26580
rect 25590 26568 25596 26580
rect 25551 26540 25596 26568
rect 25590 26528 25596 26540
rect 25648 26528 25654 26580
rect 25958 26568 25964 26580
rect 25919 26540 25964 26568
rect 25958 26528 25964 26540
rect 26016 26528 26022 26580
rect 26786 26568 26792 26580
rect 26747 26540 26792 26568
rect 26786 26528 26792 26540
rect 26844 26528 26850 26580
rect 28626 26528 28632 26580
rect 28684 26568 28690 26580
rect 28721 26571 28779 26577
rect 28721 26568 28733 26571
rect 28684 26540 28733 26568
rect 28684 26528 28690 26540
rect 28721 26537 28733 26540
rect 28767 26537 28779 26571
rect 40402 26568 40408 26580
rect 28721 26531 28779 26537
rect 31726 26540 38424 26568
rect 40363 26540 40408 26568
rect 31726 26500 31754 26540
rect 22066 26472 31754 26500
rect 8202 26432 8208 26444
rect 8163 26404 8208 26432
rect 8202 26392 8208 26404
rect 8260 26392 8266 26444
rect 16945 26435 17003 26441
rect 16945 26401 16957 26435
rect 16991 26432 17003 26435
rect 17034 26432 17040 26444
rect 16991 26404 17040 26432
rect 16991 26401 17003 26404
rect 16945 26395 17003 26401
rect 17034 26392 17040 26404
rect 17092 26392 17098 26444
rect 7469 26367 7527 26373
rect 7469 26333 7481 26367
rect 7515 26364 7527 26367
rect 7926 26364 7932 26376
rect 7515 26336 7932 26364
rect 7515 26333 7527 26336
rect 7469 26327 7527 26333
rect 7926 26324 7932 26336
rect 7984 26324 7990 26376
rect 16666 26364 16672 26376
rect 16627 26336 16672 26364
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 17310 26256 17316 26308
rect 17368 26296 17374 26308
rect 22066 26296 22094 26472
rect 33410 26460 33416 26512
rect 33468 26500 33474 26512
rect 33686 26500 33692 26512
rect 33468 26472 33692 26500
rect 33468 26460 33474 26472
rect 33686 26460 33692 26472
rect 33744 26460 33750 26512
rect 35069 26503 35127 26509
rect 35069 26469 35081 26503
rect 35115 26500 35127 26503
rect 35618 26500 35624 26512
rect 35115 26472 35624 26500
rect 35115 26469 35127 26472
rect 35069 26463 35127 26469
rect 35618 26460 35624 26472
rect 35676 26460 35682 26512
rect 35989 26503 36047 26509
rect 35989 26469 36001 26503
rect 36035 26500 36047 26503
rect 36262 26500 36268 26512
rect 36035 26472 36268 26500
rect 36035 26469 36047 26472
rect 35989 26463 36047 26469
rect 36262 26460 36268 26472
rect 36320 26460 36326 26512
rect 37734 26460 37740 26512
rect 37792 26500 37798 26512
rect 37829 26503 37887 26509
rect 37829 26500 37841 26503
rect 37792 26472 37841 26500
rect 37792 26460 37798 26472
rect 37829 26469 37841 26472
rect 37875 26469 37887 26503
rect 38286 26500 38292 26512
rect 38247 26472 38292 26500
rect 37829 26463 37887 26469
rect 38286 26460 38292 26472
rect 38344 26460 38350 26512
rect 38396 26500 38424 26540
rect 40402 26528 40408 26540
rect 40460 26528 40466 26580
rect 40770 26568 40776 26580
rect 40731 26540 40776 26568
rect 40770 26528 40776 26540
rect 40828 26528 40834 26580
rect 45370 26568 45376 26580
rect 41386 26540 45376 26568
rect 41386 26500 41414 26540
rect 45370 26528 45376 26540
rect 45428 26528 45434 26580
rect 45554 26528 45560 26580
rect 45612 26568 45618 26580
rect 45649 26571 45707 26577
rect 45649 26568 45661 26571
rect 45612 26540 45661 26568
rect 45612 26528 45618 26540
rect 45649 26537 45661 26540
rect 45695 26537 45707 26571
rect 45649 26531 45707 26537
rect 45922 26528 45928 26580
rect 45980 26568 45986 26580
rect 45980 26540 47072 26568
rect 45980 26528 45986 26540
rect 45830 26500 45836 26512
rect 38396 26472 41414 26500
rect 43272 26472 45836 26500
rect 23198 26432 23204 26444
rect 23111 26404 23204 26432
rect 23198 26392 23204 26404
rect 23256 26432 23262 26444
rect 25222 26432 25228 26444
rect 23256 26404 25228 26432
rect 23256 26392 23262 26404
rect 25222 26392 25228 26404
rect 25280 26392 25286 26444
rect 25958 26392 25964 26444
rect 26016 26432 26022 26444
rect 28350 26432 28356 26444
rect 26016 26404 26740 26432
rect 28311 26404 28356 26432
rect 26016 26392 26022 26404
rect 23014 26364 23020 26376
rect 22975 26336 23020 26364
rect 23014 26324 23020 26336
rect 23072 26364 23078 26376
rect 25774 26364 25780 26376
rect 23072 26336 25780 26364
rect 23072 26324 23078 26336
rect 25774 26324 25780 26336
rect 25832 26324 25838 26376
rect 26053 26367 26111 26373
rect 26053 26333 26065 26367
rect 26099 26364 26111 26367
rect 26234 26364 26240 26376
rect 26099 26336 26240 26364
rect 26099 26333 26111 26336
rect 26053 26327 26111 26333
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 26712 26373 26740 26404
rect 28350 26392 28356 26404
rect 28408 26392 28414 26444
rect 34698 26432 34704 26444
rect 34659 26404 34704 26432
rect 34698 26392 34704 26404
rect 34756 26392 34762 26444
rect 37642 26392 37648 26444
rect 37700 26432 37706 26444
rect 40865 26435 40923 26441
rect 37700 26404 38424 26432
rect 37700 26392 37706 26404
rect 26697 26367 26755 26373
rect 26697 26333 26709 26367
rect 26743 26333 26755 26367
rect 26697 26327 26755 26333
rect 28445 26367 28503 26373
rect 28445 26333 28457 26367
rect 28491 26364 28503 26367
rect 29638 26364 29644 26376
rect 28491 26336 29644 26364
rect 28491 26333 28503 26336
rect 28445 26327 28503 26333
rect 29638 26324 29644 26336
rect 29696 26324 29702 26376
rect 32306 26364 32312 26376
rect 32219 26336 32312 26364
rect 32306 26324 32312 26336
rect 32364 26364 32370 26376
rect 32950 26364 32956 26376
rect 32364 26336 32956 26364
rect 32364 26324 32370 26336
rect 32950 26324 32956 26336
rect 33008 26324 33014 26376
rect 34422 26324 34428 26376
rect 34480 26364 34486 26376
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34480 26336 34897 26364
rect 34480 26324 34486 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 36449 26367 36507 26373
rect 36449 26333 36461 26367
rect 36495 26364 36507 26367
rect 37826 26364 37832 26376
rect 36495 26336 37832 26364
rect 36495 26333 36507 26336
rect 36449 26327 36507 26333
rect 37826 26324 37832 26336
rect 37884 26324 37890 26376
rect 17368 26268 22094 26296
rect 32576 26299 32634 26305
rect 17368 26256 17374 26268
rect 32576 26265 32588 26299
rect 32622 26296 32634 26299
rect 32858 26296 32864 26308
rect 32622 26268 32864 26296
rect 32622 26265 32634 26268
rect 32576 26259 32634 26265
rect 32858 26256 32864 26268
rect 32916 26256 32922 26308
rect 35805 26299 35863 26305
rect 35805 26265 35817 26299
rect 35851 26296 35863 26299
rect 36716 26299 36774 26305
rect 35851 26268 36492 26296
rect 35851 26265 35863 26268
rect 35805 26259 35863 26265
rect 36464 26240 36492 26268
rect 36716 26265 36728 26299
rect 36762 26296 36774 26299
rect 36998 26296 37004 26308
rect 36762 26268 37004 26296
rect 36762 26265 36774 26268
rect 36716 26259 36774 26265
rect 36998 26256 37004 26268
rect 37056 26256 37062 26308
rect 37734 26256 37740 26308
rect 37792 26296 37798 26308
rect 37792 26268 38056 26296
rect 37792 26256 37798 26268
rect 28166 26188 28172 26240
rect 28224 26228 28230 26240
rect 29454 26228 29460 26240
rect 28224 26200 29460 26228
rect 28224 26188 28230 26200
rect 29454 26188 29460 26200
rect 29512 26188 29518 26240
rect 29730 26188 29736 26240
rect 29788 26228 29794 26240
rect 33134 26228 33140 26240
rect 29788 26200 33140 26228
rect 29788 26188 29794 26200
rect 33134 26188 33140 26200
rect 33192 26188 33198 26240
rect 36446 26188 36452 26240
rect 36504 26188 36510 26240
rect 38028 26228 38056 26268
rect 38102 26256 38108 26308
rect 38160 26296 38166 26308
rect 38289 26299 38347 26305
rect 38289 26296 38301 26299
rect 38160 26268 38301 26296
rect 38160 26256 38166 26268
rect 38289 26265 38301 26268
rect 38335 26265 38347 26299
rect 38396 26296 38424 26404
rect 40865 26401 40877 26435
rect 40911 26432 40923 26435
rect 41230 26432 41236 26444
rect 40911 26404 41236 26432
rect 40911 26401 40923 26404
rect 40865 26395 40923 26401
rect 41230 26392 41236 26404
rect 41288 26392 41294 26444
rect 43272 26432 43300 26472
rect 45830 26460 45836 26472
rect 45888 26500 45894 26512
rect 46934 26500 46940 26512
rect 45888 26472 46940 26500
rect 45888 26460 45894 26472
rect 46934 26460 46940 26472
rect 46992 26460 46998 26512
rect 41386 26404 43300 26432
rect 43349 26435 43407 26441
rect 38562 26324 38568 26376
rect 38620 26364 38626 26376
rect 38620 26336 38665 26364
rect 38620 26324 38626 26336
rect 39942 26324 39948 26376
rect 40000 26364 40006 26376
rect 40218 26364 40224 26376
rect 40000 26336 40224 26364
rect 40000 26324 40006 26336
rect 40218 26324 40224 26336
rect 40276 26324 40282 26376
rect 40586 26364 40592 26376
rect 40547 26336 40592 26364
rect 40586 26324 40592 26336
rect 40644 26324 40650 26376
rect 41386 26296 41414 26404
rect 43349 26401 43361 26435
rect 43395 26432 43407 26435
rect 43806 26432 43812 26444
rect 43395 26404 43812 26432
rect 43395 26401 43407 26404
rect 43349 26395 43407 26401
rect 43806 26392 43812 26404
rect 43864 26432 43870 26444
rect 45646 26432 45652 26444
rect 43864 26404 45652 26432
rect 43864 26392 43870 26404
rect 45646 26392 45652 26404
rect 45704 26392 45710 26444
rect 46290 26432 46296 26444
rect 46251 26404 46296 26432
rect 46290 26392 46296 26404
rect 46348 26392 46354 26444
rect 47044 26441 47072 26540
rect 47029 26435 47087 26441
rect 47029 26401 47041 26435
rect 47075 26401 47087 26435
rect 47029 26395 47087 26401
rect 45002 26364 45008 26376
rect 44963 26336 45008 26364
rect 45002 26324 45008 26336
rect 45060 26324 45066 26376
rect 45278 26364 45284 26376
rect 45239 26336 45284 26364
rect 45278 26324 45284 26336
rect 45336 26324 45342 26376
rect 45373 26367 45431 26373
rect 45373 26333 45385 26367
rect 45419 26364 45431 26367
rect 45738 26364 45744 26376
rect 45419 26336 45744 26364
rect 45419 26333 45431 26336
rect 45373 26327 45431 26333
rect 45738 26324 45744 26336
rect 45796 26324 45802 26376
rect 45922 26324 45928 26376
rect 45980 26364 45986 26376
rect 46109 26367 46167 26373
rect 46109 26364 46121 26367
rect 45980 26336 46121 26364
rect 45980 26324 45986 26336
rect 46109 26333 46121 26336
rect 46155 26333 46167 26367
rect 46109 26327 46167 26333
rect 41598 26296 41604 26308
rect 38396 26268 41414 26296
rect 41559 26268 41604 26296
rect 38289 26259 38347 26265
rect 41598 26256 41604 26268
rect 41656 26256 41662 26308
rect 44726 26256 44732 26308
rect 44784 26296 44790 26308
rect 45490 26299 45548 26305
rect 45490 26296 45502 26299
rect 44784 26268 45502 26296
rect 44784 26256 44790 26268
rect 45490 26265 45502 26268
rect 45536 26265 45548 26299
rect 45490 26259 45548 26265
rect 38473 26231 38531 26237
rect 38473 26228 38485 26231
rect 38028 26200 38485 26228
rect 38473 26197 38485 26200
rect 38519 26197 38531 26231
rect 38473 26191 38531 26197
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 26234 26024 26240 26036
rect 26195 25996 26240 26024
rect 26234 25984 26240 25996
rect 26292 25984 26298 26036
rect 27062 26024 27068 26036
rect 27023 25996 27068 26024
rect 27062 25984 27068 25996
rect 27120 26024 27126 26036
rect 27522 26024 27528 26036
rect 27120 25996 27528 26024
rect 27120 25984 27126 25996
rect 27522 25984 27528 25996
rect 27580 25984 27586 26036
rect 28442 25984 28448 26036
rect 28500 26024 28506 26036
rect 28629 26027 28687 26033
rect 28629 26024 28641 26027
rect 28500 25996 28641 26024
rect 28500 25984 28506 25996
rect 28629 25993 28641 25996
rect 28675 25993 28687 26027
rect 29917 26027 29975 26033
rect 28629 25987 28687 25993
rect 28828 25996 29868 26024
rect 8570 25916 8576 25968
rect 8628 25956 8634 25968
rect 28828 25956 28856 25996
rect 29549 25959 29607 25965
rect 29549 25956 29561 25959
rect 8628 25928 28856 25956
rect 28920 25928 29561 25956
rect 8628 25916 8634 25928
rect 7834 25848 7840 25900
rect 7892 25888 7898 25900
rect 8021 25891 8079 25897
rect 8021 25888 8033 25891
rect 7892 25860 8033 25888
rect 7892 25848 7898 25860
rect 8021 25857 8033 25860
rect 8067 25888 8079 25891
rect 9217 25891 9275 25897
rect 9217 25888 9229 25891
rect 8067 25860 9229 25888
rect 8067 25857 8079 25860
rect 8021 25851 8079 25857
rect 9217 25857 9229 25860
rect 9263 25857 9275 25891
rect 9217 25851 9275 25857
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25888 22247 25891
rect 23474 25888 23480 25900
rect 22235 25860 23480 25888
rect 22235 25857 22247 25860
rect 22189 25851 22247 25857
rect 23474 25848 23480 25860
rect 23532 25848 23538 25900
rect 25124 25891 25182 25897
rect 25124 25857 25136 25891
rect 25170 25888 25182 25891
rect 25498 25888 25504 25900
rect 25170 25860 25504 25888
rect 25170 25857 25182 25860
rect 25124 25851 25182 25857
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 26234 25848 26240 25900
rect 26292 25888 26298 25900
rect 26973 25891 27031 25897
rect 26973 25888 26985 25891
rect 26292 25860 26985 25888
rect 26292 25848 26298 25860
rect 26973 25857 26985 25860
rect 27019 25857 27031 25891
rect 27982 25888 27988 25900
rect 27943 25860 27988 25888
rect 26973 25851 27031 25857
rect 27982 25848 27988 25860
rect 28040 25848 28046 25900
rect 28166 25888 28172 25900
rect 28127 25860 28172 25888
rect 28166 25848 28172 25860
rect 28224 25848 28230 25900
rect 28350 25848 28356 25900
rect 28408 25888 28414 25900
rect 28813 25891 28871 25897
rect 28813 25888 28825 25891
rect 28408 25860 28825 25888
rect 28408 25848 28414 25860
rect 28813 25857 28825 25860
rect 28859 25857 28871 25891
rect 28813 25851 28871 25857
rect 28920 25832 28948 25928
rect 29549 25925 29561 25928
rect 29595 25925 29607 25959
rect 29749 25959 29807 25965
rect 29749 25956 29761 25959
rect 29549 25919 29607 25925
rect 29656 25928 29761 25956
rect 28994 25848 29000 25900
rect 29052 25888 29058 25900
rect 29656 25888 29684 25928
rect 29749 25925 29761 25928
rect 29795 25925 29807 25959
rect 29749 25919 29807 25925
rect 29052 25860 29684 25888
rect 29052 25848 29058 25860
rect 8570 25820 8576 25832
rect 8531 25792 8576 25820
rect 8570 25780 8576 25792
rect 8628 25780 8634 25832
rect 9490 25820 9496 25832
rect 9451 25792 9496 25820
rect 9490 25780 9496 25792
rect 9548 25780 9554 25832
rect 22281 25823 22339 25829
rect 22281 25789 22293 25823
rect 22327 25820 22339 25823
rect 23198 25820 23204 25832
rect 22327 25792 23204 25820
rect 22327 25789 22339 25792
rect 22281 25783 22339 25789
rect 23198 25780 23204 25792
rect 23256 25780 23262 25832
rect 24854 25820 24860 25832
rect 24815 25792 24860 25820
rect 24854 25780 24860 25792
rect 24912 25780 24918 25832
rect 28902 25780 28908 25832
rect 28960 25780 28966 25832
rect 29086 25820 29092 25832
rect 29047 25792 29092 25820
rect 29086 25780 29092 25792
rect 29144 25780 29150 25832
rect 3050 25712 3056 25764
rect 3108 25752 3114 25764
rect 9508 25752 9536 25780
rect 3108 25724 9536 25752
rect 3108 25712 3114 25724
rect 28718 25712 28724 25764
rect 28776 25752 28782 25764
rect 29840 25752 29868 25996
rect 29917 25993 29929 26027
rect 29963 26024 29975 26027
rect 33781 26027 33839 26033
rect 29963 25996 30788 26024
rect 29963 25993 29975 25996
rect 29917 25987 29975 25993
rect 30558 25888 30564 25900
rect 30519 25860 30564 25888
rect 30558 25848 30564 25860
rect 30616 25848 30622 25900
rect 30760 25897 30788 25996
rect 33781 25993 33793 26027
rect 33827 26024 33839 26027
rect 34422 26024 34428 26036
rect 33827 25996 34428 26024
rect 33827 25993 33839 25996
rect 33781 25987 33839 25993
rect 34422 25984 34428 25996
rect 34480 25984 34486 26036
rect 39850 25984 39856 26036
rect 39908 26024 39914 26036
rect 40313 26027 40371 26033
rect 40313 26024 40325 26027
rect 39908 25996 40325 26024
rect 39908 25984 39914 25996
rect 40313 25993 40325 25996
rect 40359 25993 40371 26027
rect 40313 25987 40371 25993
rect 32677 25959 32735 25965
rect 32677 25925 32689 25959
rect 32723 25956 32735 25959
rect 33410 25956 33416 25968
rect 32723 25928 33416 25956
rect 32723 25925 32735 25928
rect 32677 25919 32735 25925
rect 33410 25916 33416 25928
rect 33468 25916 33474 25968
rect 33613 25959 33671 25965
rect 33613 25956 33625 25959
rect 33520 25928 33625 25956
rect 30745 25891 30803 25897
rect 30745 25857 30757 25891
rect 30791 25857 30803 25891
rect 31110 25888 31116 25900
rect 31071 25860 31116 25888
rect 30745 25851 30803 25857
rect 31110 25848 31116 25860
rect 31168 25848 31174 25900
rect 32861 25891 32919 25897
rect 32861 25857 32873 25891
rect 32907 25857 32919 25891
rect 32861 25851 32919 25857
rect 32953 25891 33011 25897
rect 32953 25857 32965 25891
rect 32999 25888 33011 25891
rect 33134 25888 33140 25900
rect 32999 25860 33140 25888
rect 32999 25857 33011 25860
rect 32953 25851 33011 25857
rect 29914 25780 29920 25832
rect 29972 25820 29978 25832
rect 30837 25823 30895 25829
rect 30837 25820 30849 25823
rect 29972 25792 30849 25820
rect 29972 25780 29978 25792
rect 30837 25789 30849 25792
rect 30883 25789 30895 25823
rect 30837 25783 30895 25789
rect 30929 25823 30987 25829
rect 30929 25789 30941 25823
rect 30975 25820 30987 25823
rect 32398 25820 32404 25832
rect 30975 25792 32404 25820
rect 30975 25789 30987 25792
rect 30929 25783 30987 25789
rect 32398 25780 32404 25792
rect 32456 25780 32462 25832
rect 32876 25820 32904 25851
rect 33134 25848 33140 25860
rect 33192 25888 33198 25900
rect 33520 25888 33548 25928
rect 33613 25925 33625 25928
rect 33659 25925 33671 25959
rect 41874 25956 41880 25968
rect 33613 25919 33671 25925
rect 33704 25928 41880 25956
rect 33192 25860 33548 25888
rect 33192 25848 33198 25860
rect 33594 25820 33600 25832
rect 32876 25792 33600 25820
rect 33594 25780 33600 25792
rect 33652 25780 33658 25832
rect 32674 25752 32680 25764
rect 28776 25724 29776 25752
rect 29840 25724 31754 25752
rect 32635 25724 32680 25752
rect 28776 25712 28782 25724
rect 22462 25684 22468 25696
rect 22423 25656 22468 25684
rect 22462 25644 22468 25656
rect 22520 25644 22526 25696
rect 28077 25687 28135 25693
rect 28077 25653 28089 25687
rect 28123 25684 28135 25687
rect 28902 25684 28908 25696
rect 28123 25656 28908 25684
rect 28123 25653 28135 25656
rect 28077 25647 28135 25653
rect 28902 25644 28908 25656
rect 28960 25644 28966 25696
rect 28997 25687 29055 25693
rect 28997 25653 29009 25687
rect 29043 25684 29055 25687
rect 29454 25684 29460 25696
rect 29043 25656 29460 25684
rect 29043 25653 29055 25656
rect 28997 25647 29055 25653
rect 29454 25644 29460 25656
rect 29512 25644 29518 25696
rect 29748 25693 29776 25724
rect 29733 25687 29791 25693
rect 29733 25653 29745 25687
rect 29779 25653 29791 25687
rect 31294 25684 31300 25696
rect 31255 25656 31300 25684
rect 29733 25647 29791 25653
rect 31294 25644 31300 25656
rect 31352 25644 31358 25696
rect 31726 25684 31754 25724
rect 32674 25712 32680 25724
rect 32732 25712 32738 25764
rect 33704 25752 33732 25928
rect 41874 25916 41880 25928
rect 41932 25916 41938 25968
rect 44266 25916 44272 25968
rect 44324 25956 44330 25968
rect 45833 25959 45891 25965
rect 45833 25956 45845 25959
rect 44324 25928 45845 25956
rect 44324 25916 44330 25928
rect 45833 25925 45845 25928
rect 45879 25925 45891 25959
rect 45833 25919 45891 25925
rect 36446 25888 36452 25900
rect 36407 25860 36452 25888
rect 36446 25848 36452 25860
rect 36504 25848 36510 25900
rect 39022 25888 39028 25900
rect 38983 25860 39028 25888
rect 39022 25848 39028 25860
rect 39080 25888 39086 25900
rect 41598 25888 41604 25900
rect 39080 25860 41604 25888
rect 39080 25848 39086 25860
rect 41598 25848 41604 25860
rect 41656 25848 41662 25900
rect 43625 25891 43683 25897
rect 43625 25857 43637 25891
rect 43671 25888 43683 25891
rect 45002 25888 45008 25900
rect 43671 25860 45008 25888
rect 43671 25857 43683 25860
rect 43625 25851 43683 25857
rect 44545 25823 44603 25829
rect 44545 25820 44557 25823
rect 44008 25792 44557 25820
rect 44008 25761 44036 25792
rect 44545 25789 44557 25792
rect 44591 25820 44603 25823
rect 44726 25820 44732 25832
rect 44591 25792 44732 25820
rect 44591 25789 44603 25792
rect 44545 25783 44603 25789
rect 44726 25780 44732 25792
rect 44784 25780 44790 25832
rect 44836 25761 44864 25860
rect 45002 25848 45008 25860
rect 45060 25848 45066 25900
rect 45278 25848 45284 25900
rect 45336 25888 45342 25900
rect 45465 25891 45523 25897
rect 45465 25888 45477 25891
rect 45336 25860 45477 25888
rect 45336 25848 45342 25860
rect 45465 25857 45477 25860
rect 45511 25857 45523 25891
rect 45465 25851 45523 25857
rect 45649 25891 45707 25897
rect 45649 25857 45661 25891
rect 45695 25888 45707 25891
rect 45738 25888 45744 25900
rect 45695 25860 45744 25888
rect 45695 25857 45707 25860
rect 45649 25851 45707 25857
rect 45480 25820 45508 25851
rect 45738 25848 45744 25860
rect 45796 25888 45802 25900
rect 46293 25891 46351 25897
rect 46293 25888 46305 25891
rect 45796 25860 46305 25888
rect 45796 25848 45802 25860
rect 46293 25857 46305 25860
rect 46339 25857 46351 25891
rect 46293 25851 46351 25857
rect 46477 25891 46535 25897
rect 46477 25857 46489 25891
rect 46523 25857 46535 25891
rect 46477 25851 46535 25857
rect 46492 25820 46520 25851
rect 46934 25848 46940 25900
rect 46992 25888 46998 25900
rect 47581 25891 47639 25897
rect 47581 25888 47593 25891
rect 46992 25860 47593 25888
rect 46992 25848 46998 25860
rect 47581 25857 47593 25860
rect 47627 25857 47639 25891
rect 47581 25851 47639 25857
rect 45480 25792 46520 25820
rect 33520 25724 33732 25752
rect 43993 25755 44051 25761
rect 33520 25684 33548 25724
rect 43993 25721 44005 25755
rect 44039 25721 44051 25755
rect 43993 25715 44051 25721
rect 44821 25755 44879 25761
rect 44821 25721 44833 25755
rect 44867 25721 44879 25755
rect 46293 25755 46351 25761
rect 46293 25752 46305 25755
rect 44821 25715 44879 25721
rect 45480 25724 46305 25752
rect 45480 25696 45508 25724
rect 46293 25721 46305 25724
rect 46339 25721 46351 25755
rect 46293 25715 46351 25721
rect 31726 25656 33548 25684
rect 33594 25644 33600 25696
rect 33652 25684 33658 25696
rect 33870 25684 33876 25696
rect 33652 25656 33876 25684
rect 33652 25644 33658 25656
rect 33870 25644 33876 25656
rect 33928 25644 33934 25696
rect 36538 25684 36544 25696
rect 36499 25656 36544 25684
rect 36538 25644 36544 25656
rect 36596 25684 36602 25696
rect 38930 25684 38936 25696
rect 36596 25656 38936 25684
rect 36596 25644 36602 25656
rect 38930 25644 38936 25656
rect 38988 25684 38994 25696
rect 39942 25684 39948 25696
rect 38988 25656 39948 25684
rect 38988 25644 38994 25656
rect 39942 25644 39948 25656
rect 40000 25644 40006 25696
rect 44085 25687 44143 25693
rect 44085 25653 44097 25687
rect 44131 25684 44143 25687
rect 44358 25684 44364 25696
rect 44131 25656 44364 25684
rect 44131 25653 44143 25656
rect 44085 25647 44143 25653
rect 44358 25644 44364 25656
rect 44416 25644 44422 25696
rect 45005 25687 45063 25693
rect 45005 25653 45017 25687
rect 45051 25684 45063 25687
rect 45370 25684 45376 25696
rect 45051 25656 45376 25684
rect 45051 25653 45063 25656
rect 45005 25647 45063 25653
rect 45370 25644 45376 25656
rect 45428 25644 45434 25696
rect 45462 25644 45468 25696
rect 45520 25644 45526 25696
rect 46474 25644 46480 25696
rect 46532 25684 46538 25696
rect 47673 25687 47731 25693
rect 47673 25684 47685 25687
rect 46532 25656 47685 25684
rect 46532 25644 46538 25656
rect 47673 25653 47685 25656
rect 47719 25653 47731 25687
rect 47673 25647 47731 25653
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 25498 25480 25504 25492
rect 25459 25452 25504 25480
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 29086 25480 29092 25492
rect 27908 25452 29092 25480
rect 25409 25415 25467 25421
rect 25409 25381 25421 25415
rect 25455 25412 25467 25415
rect 26053 25415 26111 25421
rect 26053 25412 26065 25415
rect 25455 25384 26065 25412
rect 25455 25381 25467 25384
rect 25409 25375 25467 25381
rect 26053 25381 26065 25384
rect 26099 25381 26111 25415
rect 26053 25375 26111 25381
rect 18782 25344 18788 25356
rect 6886 25316 18788 25344
rect 2130 25276 2136 25288
rect 2091 25248 2136 25276
rect 2130 25236 2136 25248
rect 2188 25236 2194 25288
rect 2593 25279 2651 25285
rect 2593 25245 2605 25279
rect 2639 25276 2651 25279
rect 6886 25276 6914 25316
rect 18782 25304 18788 25316
rect 18840 25304 18846 25356
rect 27614 25344 27620 25356
rect 22020 25316 22692 25344
rect 7834 25276 7840 25288
rect 2639 25248 6914 25276
rect 7795 25248 7840 25276
rect 2639 25245 2651 25248
rect 2593 25239 2651 25245
rect 7834 25236 7840 25248
rect 7892 25236 7898 25288
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25276 8171 25279
rect 12526 25276 12532 25288
rect 8159 25248 12532 25276
rect 8159 25245 8171 25248
rect 8113 25239 8171 25245
rect 12526 25236 12532 25248
rect 12584 25236 12590 25288
rect 22020 25285 22048 25316
rect 22664 25288 22692 25316
rect 23308 25316 27620 25344
rect 21821 25279 21879 25285
rect 21821 25245 21833 25279
rect 21867 25245 21879 25279
rect 21821 25239 21879 25245
rect 22005 25279 22063 25285
rect 22005 25245 22017 25279
rect 22051 25245 22063 25279
rect 22462 25276 22468 25288
rect 22423 25248 22468 25276
rect 22005 25239 22063 25245
rect 21836 25208 21864 25239
rect 22462 25236 22468 25248
rect 22520 25236 22526 25288
rect 22646 25276 22652 25288
rect 22607 25248 22652 25276
rect 22646 25236 22652 25248
rect 22704 25236 22710 25288
rect 23106 25236 23112 25288
rect 23164 25276 23170 25288
rect 23308 25285 23336 25316
rect 23293 25279 23351 25285
rect 23293 25276 23305 25279
rect 23164 25248 23305 25276
rect 23164 25236 23170 25248
rect 23293 25245 23305 25248
rect 23339 25245 23351 25279
rect 23474 25276 23480 25288
rect 23435 25248 23480 25276
rect 23293 25239 23351 25245
rect 23474 25236 23480 25248
rect 23532 25236 23538 25288
rect 25130 25276 25136 25288
rect 25091 25248 25136 25276
rect 25130 25236 25136 25248
rect 25188 25236 25194 25288
rect 25314 25276 25320 25288
rect 25275 25248 25320 25276
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 26068 25285 26096 25316
rect 27614 25304 27620 25316
rect 27672 25304 27678 25356
rect 25501 25279 25559 25285
rect 25501 25245 25513 25279
rect 25547 25245 25559 25279
rect 25501 25239 25559 25245
rect 26053 25279 26111 25285
rect 26053 25245 26065 25279
rect 26099 25245 26111 25279
rect 26234 25276 26240 25288
rect 26195 25248 26240 25276
rect 26053 25239 26111 25245
rect 22480 25208 22508 25236
rect 21836 25180 22508 25208
rect 25516 25208 25544 25239
rect 26234 25236 26240 25248
rect 26292 25236 26298 25288
rect 27908 25285 27936 25452
rect 29086 25440 29092 25452
rect 29144 25480 29150 25492
rect 31110 25480 31116 25492
rect 29144 25452 31116 25480
rect 29144 25440 29150 25452
rect 31110 25440 31116 25452
rect 31168 25480 31174 25492
rect 32125 25483 32183 25489
rect 32125 25480 32137 25483
rect 31168 25452 32137 25480
rect 31168 25440 31174 25452
rect 32125 25449 32137 25452
rect 32171 25449 32183 25483
rect 32125 25443 32183 25449
rect 33318 25440 33324 25492
rect 33376 25480 33382 25492
rect 36538 25480 36544 25492
rect 33376 25452 36544 25480
rect 33376 25440 33382 25452
rect 36538 25440 36544 25452
rect 36596 25440 36602 25492
rect 40310 25440 40316 25492
rect 40368 25480 40374 25492
rect 40405 25483 40463 25489
rect 40405 25480 40417 25483
rect 40368 25452 40417 25480
rect 40368 25440 40374 25452
rect 40405 25449 40417 25452
rect 40451 25449 40463 25483
rect 44358 25480 44364 25492
rect 44319 25452 44364 25480
rect 40405 25443 40463 25449
rect 28718 25372 28724 25424
rect 28776 25372 28782 25424
rect 29638 25412 29644 25424
rect 29599 25384 29644 25412
rect 29638 25372 29644 25384
rect 29696 25412 29702 25424
rect 30374 25412 30380 25424
rect 29696 25384 30380 25412
rect 29696 25372 29702 25384
rect 30374 25372 30380 25384
rect 30432 25372 30438 25424
rect 35802 25412 35808 25424
rect 35763 25384 35808 25412
rect 35802 25372 35808 25384
rect 35860 25372 35866 25424
rect 28736 25344 28764 25372
rect 40420 25344 40448 25443
rect 44358 25440 44364 25452
rect 44416 25440 44422 25492
rect 45278 25412 45284 25424
rect 44376 25384 45284 25412
rect 41598 25344 41604 25356
rect 28736 25316 29040 25344
rect 40420 25316 41604 25344
rect 27893 25279 27951 25285
rect 27893 25245 27905 25279
rect 27939 25245 27951 25279
rect 27893 25239 27951 25245
rect 28534 25236 28540 25288
rect 28592 25276 28598 25288
rect 28718 25276 28724 25288
rect 28592 25248 28724 25276
rect 28592 25236 28598 25248
rect 28718 25236 28724 25248
rect 28776 25236 28782 25288
rect 28902 25276 28908 25288
rect 28863 25248 28908 25276
rect 28902 25236 28908 25248
rect 28960 25236 28966 25288
rect 29012 25285 29040 25316
rect 41598 25304 41604 25316
rect 41656 25304 41662 25356
rect 44266 25344 44272 25356
rect 44100 25316 44272 25344
rect 28997 25279 29055 25285
rect 28997 25245 29009 25279
rect 29043 25245 29055 25279
rect 28997 25239 29055 25245
rect 29454 25236 29460 25288
rect 29512 25276 29518 25288
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 29512 25248 29561 25276
rect 29512 25236 29518 25248
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 30745 25279 30803 25285
rect 30745 25245 30757 25279
rect 30791 25276 30803 25279
rect 32306 25276 32312 25288
rect 30791 25248 32312 25276
rect 30791 25245 30803 25248
rect 30745 25239 30803 25245
rect 32306 25236 32312 25248
rect 32364 25236 32370 25288
rect 35805 25279 35863 25285
rect 35805 25245 35817 25279
rect 35851 25276 35863 25279
rect 35894 25276 35900 25288
rect 35851 25248 35900 25276
rect 35851 25245 35863 25248
rect 35805 25239 35863 25245
rect 35894 25236 35900 25248
rect 35952 25236 35958 25288
rect 35986 25236 35992 25288
rect 36044 25276 36050 25288
rect 40954 25276 40960 25288
rect 36044 25248 36089 25276
rect 40915 25248 40960 25276
rect 36044 25236 36050 25248
rect 40954 25236 40960 25248
rect 41012 25236 41018 25288
rect 44100 25285 44128 25316
rect 44266 25304 44272 25316
rect 44324 25304 44330 25356
rect 44085 25279 44143 25285
rect 44085 25245 44097 25279
rect 44131 25245 44143 25279
rect 44085 25239 44143 25245
rect 44174 25236 44180 25288
rect 44232 25276 44238 25288
rect 44376 25276 44404 25384
rect 45278 25372 45284 25384
rect 45336 25412 45342 25424
rect 45462 25412 45468 25424
rect 45336 25384 45468 25412
rect 45336 25372 45342 25384
rect 45462 25372 45468 25384
rect 45520 25372 45526 25424
rect 44542 25344 44548 25356
rect 44455 25316 44548 25344
rect 44468 25285 44496 25316
rect 44542 25304 44548 25316
rect 44600 25344 44606 25356
rect 44600 25316 45416 25344
rect 44600 25304 44606 25316
rect 45388 25288 45416 25316
rect 44232 25248 44404 25276
rect 44453 25279 44511 25285
rect 44232 25236 44238 25248
rect 44453 25245 44465 25279
rect 44499 25245 44511 25279
rect 44453 25239 44511 25245
rect 45189 25279 45247 25285
rect 45189 25245 45201 25279
rect 45235 25245 45247 25279
rect 45370 25276 45376 25288
rect 45331 25248 45376 25276
rect 45189 25239 45247 25245
rect 29730 25208 29736 25220
rect 25516 25180 29736 25208
rect 29730 25168 29736 25180
rect 29788 25168 29794 25220
rect 31012 25211 31070 25217
rect 31012 25177 31024 25211
rect 31058 25208 31070 25211
rect 31294 25208 31300 25220
rect 31058 25180 31300 25208
rect 31058 25177 31070 25180
rect 31012 25171 31070 25177
rect 31294 25168 31300 25180
rect 31352 25168 31358 25220
rect 36446 25168 36452 25220
rect 36504 25208 36510 25220
rect 40313 25211 40371 25217
rect 40313 25208 40325 25211
rect 36504 25180 40325 25208
rect 36504 25168 36510 25180
rect 40313 25177 40325 25180
rect 40359 25208 40371 25211
rect 43438 25208 43444 25220
rect 40359 25180 43444 25208
rect 40359 25177 40371 25180
rect 40313 25171 40371 25177
rect 43438 25168 43444 25180
rect 43496 25168 43502 25220
rect 45204 25208 45232 25239
rect 45370 25236 45376 25248
rect 45428 25236 45434 25288
rect 45480 25285 45508 25372
rect 46474 25344 46480 25356
rect 46435 25316 46480 25344
rect 46474 25304 46480 25316
rect 46532 25304 46538 25356
rect 46750 25344 46756 25356
rect 46711 25316 46756 25344
rect 46750 25304 46756 25316
rect 46808 25304 46814 25356
rect 45465 25279 45523 25285
rect 45465 25245 45477 25279
rect 45511 25245 45523 25279
rect 45465 25239 45523 25245
rect 46293 25279 46351 25285
rect 46293 25245 46305 25279
rect 46339 25245 46351 25279
rect 46293 25239 46351 25245
rect 45554 25208 45560 25220
rect 45204 25180 45560 25208
rect 45554 25168 45560 25180
rect 45612 25168 45618 25220
rect 46308 25208 46336 25239
rect 47762 25208 47768 25220
rect 46308 25180 47768 25208
rect 47762 25168 47768 25180
rect 47820 25168 47826 25220
rect 2314 25100 2320 25152
rect 2372 25140 2378 25152
rect 2685 25143 2743 25149
rect 2685 25140 2697 25143
rect 2372 25112 2697 25140
rect 2372 25100 2378 25112
rect 2685 25109 2697 25112
rect 2731 25109 2743 25143
rect 2685 25103 2743 25109
rect 22005 25143 22063 25149
rect 22005 25109 22017 25143
rect 22051 25140 22063 25143
rect 22738 25140 22744 25152
rect 22051 25112 22744 25140
rect 22051 25109 22063 25112
rect 22005 25103 22063 25109
rect 22738 25100 22744 25112
rect 22796 25100 22802 25152
rect 22833 25143 22891 25149
rect 22833 25109 22845 25143
rect 22879 25140 22891 25143
rect 22922 25140 22928 25152
rect 22879 25112 22928 25140
rect 22879 25109 22891 25112
rect 22833 25103 22891 25109
rect 22922 25100 22928 25112
rect 22980 25100 22986 25152
rect 23290 25100 23296 25152
rect 23348 25140 23354 25152
rect 23385 25143 23443 25149
rect 23385 25140 23397 25143
rect 23348 25112 23397 25140
rect 23348 25100 23354 25112
rect 23385 25109 23397 25112
rect 23431 25109 23443 25143
rect 23385 25103 23443 25109
rect 27798 25100 27804 25152
rect 27856 25140 27862 25152
rect 27985 25143 28043 25149
rect 27985 25140 27997 25143
rect 27856 25112 27997 25140
rect 27856 25100 27862 25112
rect 27985 25109 27997 25112
rect 28031 25109 28043 25143
rect 27985 25103 28043 25109
rect 28537 25143 28595 25149
rect 28537 25109 28549 25143
rect 28583 25140 28595 25143
rect 28626 25140 28632 25152
rect 28583 25112 28632 25140
rect 28583 25109 28595 25112
rect 28537 25103 28595 25109
rect 28626 25100 28632 25112
rect 28684 25100 28690 25152
rect 41049 25143 41107 25149
rect 41049 25109 41061 25143
rect 41095 25140 41107 25143
rect 41414 25140 41420 25152
rect 41095 25112 41420 25140
rect 41095 25109 41107 25112
rect 41049 25103 41107 25109
rect 41414 25100 41420 25112
rect 41472 25100 41478 25152
rect 43901 25143 43959 25149
rect 43901 25109 43913 25143
rect 43947 25140 43959 25143
rect 44910 25140 44916 25152
rect 43947 25112 44916 25140
rect 43947 25109 43959 25112
rect 43901 25103 43959 25109
rect 44910 25100 44916 25112
rect 44968 25100 44974 25152
rect 45005 25143 45063 25149
rect 45005 25109 45017 25143
rect 45051 25140 45063 25143
rect 45186 25140 45192 25152
rect 45051 25112 45192 25140
rect 45051 25109 45063 25112
rect 45005 25103 45063 25109
rect 45186 25100 45192 25112
rect 45244 25100 45250 25152
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 28169 24939 28227 24945
rect 28169 24905 28181 24939
rect 28215 24936 28227 24939
rect 28718 24936 28724 24948
rect 28215 24908 28724 24936
rect 28215 24905 28227 24908
rect 28169 24899 28227 24905
rect 28718 24896 28724 24908
rect 28776 24896 28782 24948
rect 33686 24896 33692 24948
rect 33744 24936 33750 24948
rect 40954 24936 40960 24948
rect 33744 24908 40960 24936
rect 33744 24896 33750 24908
rect 40954 24896 40960 24908
rect 41012 24896 41018 24948
rect 2314 24868 2320 24880
rect 2275 24840 2320 24868
rect 2314 24828 2320 24840
rect 2372 24828 2378 24880
rect 27614 24828 27620 24880
rect 27672 24868 27678 24880
rect 38746 24868 38752 24880
rect 27672 24840 28856 24868
rect 27672 24828 27678 24840
rect 2130 24800 2136 24812
rect 2091 24772 2136 24800
rect 2130 24760 2136 24772
rect 2188 24760 2194 24812
rect 7834 24800 7840 24812
rect 7795 24772 7840 24800
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 23474 24760 23480 24812
rect 23532 24800 23538 24812
rect 24762 24800 24768 24812
rect 23532 24772 24768 24800
rect 23532 24760 23538 24772
rect 24762 24760 24768 24772
rect 24820 24760 24826 24812
rect 27798 24800 27804 24812
rect 27759 24772 27804 24800
rect 27798 24760 27804 24772
rect 27856 24760 27862 24812
rect 28626 24800 28632 24812
rect 28587 24772 28632 24800
rect 28626 24760 28632 24772
rect 28684 24760 28690 24812
rect 28828 24809 28856 24840
rect 38212 24840 38752 24868
rect 28813 24803 28871 24809
rect 28813 24769 28825 24803
rect 28859 24769 28871 24803
rect 28813 24763 28871 24769
rect 31021 24803 31079 24809
rect 31021 24769 31033 24803
rect 31067 24800 31079 24803
rect 32214 24800 32220 24812
rect 31067 24772 32220 24800
rect 31067 24769 31079 24772
rect 31021 24763 31079 24769
rect 32214 24760 32220 24772
rect 32272 24760 32278 24812
rect 35710 24760 35716 24812
rect 35768 24800 35774 24812
rect 35805 24803 35863 24809
rect 35805 24800 35817 24803
rect 35768 24772 35817 24800
rect 35768 24760 35774 24772
rect 35805 24769 35817 24772
rect 35851 24769 35863 24803
rect 35805 24763 35863 24769
rect 36449 24803 36507 24809
rect 36449 24769 36461 24803
rect 36495 24800 36507 24803
rect 37274 24800 37280 24812
rect 36495 24772 37280 24800
rect 36495 24769 36507 24772
rect 36449 24763 36507 24769
rect 37274 24760 37280 24772
rect 37332 24760 37338 24812
rect 38013 24803 38071 24809
rect 38013 24769 38025 24803
rect 38059 24800 38071 24803
rect 38212 24800 38240 24840
rect 38746 24828 38752 24840
rect 38804 24828 38810 24880
rect 44358 24868 44364 24880
rect 44284 24840 44364 24868
rect 38059 24772 38240 24800
rect 38280 24803 38338 24809
rect 38059 24769 38071 24772
rect 38013 24763 38071 24769
rect 38280 24769 38292 24803
rect 38326 24800 38338 24803
rect 39482 24800 39488 24812
rect 38326 24772 39488 24800
rect 38326 24769 38338 24772
rect 38280 24763 38338 24769
rect 39482 24760 39488 24772
rect 39540 24760 39546 24812
rect 39574 24760 39580 24812
rect 39632 24800 39638 24812
rect 39853 24803 39911 24809
rect 39853 24800 39865 24803
rect 39632 24772 39865 24800
rect 39632 24760 39638 24772
rect 39853 24769 39865 24772
rect 39899 24769 39911 24803
rect 39853 24763 39911 24769
rect 40037 24803 40095 24809
rect 40037 24769 40049 24803
rect 40083 24769 40095 24803
rect 40037 24763 40095 24769
rect 2774 24732 2780 24744
rect 2735 24704 2780 24732
rect 2774 24692 2780 24704
rect 2832 24692 2838 24744
rect 8018 24732 8024 24744
rect 7979 24704 8024 24732
rect 8018 24692 8024 24704
rect 8076 24692 8082 24744
rect 22002 24732 22008 24744
rect 21963 24704 22008 24732
rect 22002 24692 22008 24704
rect 22060 24692 22066 24744
rect 22186 24732 22192 24744
rect 22147 24704 22192 24732
rect 22186 24692 22192 24704
rect 22244 24692 22250 24744
rect 22465 24735 22523 24741
rect 22465 24701 22477 24735
rect 22511 24701 22523 24735
rect 22465 24695 22523 24701
rect 27893 24735 27951 24741
rect 27893 24701 27905 24735
rect 27939 24732 27951 24735
rect 28350 24732 28356 24744
rect 27939 24704 28356 24732
rect 27939 24701 27951 24704
rect 27893 24695 27951 24701
rect 3418 24624 3424 24676
rect 3476 24664 3482 24676
rect 22480 24664 22508 24695
rect 28350 24692 28356 24704
rect 28408 24692 28414 24744
rect 28721 24735 28779 24741
rect 28721 24701 28733 24735
rect 28767 24732 28779 24735
rect 29914 24732 29920 24744
rect 28767 24704 29920 24732
rect 28767 24701 28779 24704
rect 28721 24695 28779 24701
rect 29914 24692 29920 24704
rect 29972 24692 29978 24744
rect 33321 24735 33379 24741
rect 33321 24701 33333 24735
rect 33367 24732 33379 24735
rect 33410 24732 33416 24744
rect 33367 24704 33416 24732
rect 33367 24701 33379 24704
rect 33321 24695 33379 24701
rect 33410 24692 33416 24704
rect 33468 24692 33474 24744
rect 33597 24735 33655 24741
rect 33597 24701 33609 24735
rect 33643 24732 33655 24735
rect 33962 24732 33968 24744
rect 33643 24704 33968 24732
rect 33643 24701 33655 24704
rect 33597 24695 33655 24701
rect 33962 24692 33968 24704
rect 34020 24692 34026 24744
rect 35526 24692 35532 24744
rect 35584 24732 35590 24744
rect 35621 24735 35679 24741
rect 35621 24732 35633 24735
rect 35584 24704 35633 24732
rect 35584 24692 35590 24704
rect 35621 24701 35633 24704
rect 35667 24701 35679 24735
rect 35621 24695 35679 24701
rect 36725 24735 36783 24741
rect 36725 24701 36737 24735
rect 36771 24701 36783 24735
rect 36725 24695 36783 24701
rect 3476 24636 22508 24664
rect 3476 24624 3482 24636
rect 35894 24624 35900 24676
rect 35952 24664 35958 24676
rect 36633 24667 36691 24673
rect 36633 24664 36645 24667
rect 35952 24636 36645 24664
rect 35952 24624 35958 24636
rect 36633 24633 36645 24636
rect 36679 24633 36691 24667
rect 36743 24664 36771 24695
rect 39114 24692 39120 24744
rect 39172 24732 39178 24744
rect 40052 24732 40080 24763
rect 43254 24760 43260 24812
rect 43312 24800 43318 24812
rect 43993 24803 44051 24809
rect 43993 24800 44005 24803
rect 43312 24772 44005 24800
rect 43312 24760 43318 24772
rect 43993 24769 44005 24772
rect 44039 24769 44051 24803
rect 44174 24800 44180 24812
rect 44135 24772 44180 24800
rect 43993 24763 44051 24769
rect 44174 24760 44180 24772
rect 44232 24760 44238 24812
rect 44284 24809 44312 24840
rect 44358 24828 44364 24840
rect 44416 24828 44422 24880
rect 45554 24828 45560 24880
rect 45612 24868 45618 24880
rect 45612 24840 45692 24868
rect 45612 24828 45618 24840
rect 44269 24803 44327 24809
rect 44269 24769 44281 24803
rect 44315 24769 44327 24803
rect 44542 24800 44548 24812
rect 44503 24772 44548 24800
rect 44269 24763 44327 24769
rect 44542 24760 44548 24772
rect 44600 24760 44606 24812
rect 45278 24760 45284 24812
rect 45336 24800 45342 24812
rect 45373 24803 45431 24809
rect 45373 24800 45385 24803
rect 45336 24772 45385 24800
rect 45336 24760 45342 24772
rect 45373 24769 45385 24772
rect 45419 24769 45431 24803
rect 45373 24763 45431 24769
rect 45462 24760 45468 24812
rect 45520 24800 45526 24812
rect 45664 24809 45692 24840
rect 45649 24803 45707 24809
rect 45520 24772 45565 24800
rect 45520 24760 45526 24772
rect 45649 24769 45661 24803
rect 45695 24769 45707 24803
rect 45649 24763 45707 24769
rect 45741 24803 45799 24809
rect 45741 24769 45753 24803
rect 45787 24800 45799 24803
rect 46293 24803 46351 24809
rect 46293 24800 46305 24803
rect 45787 24772 46305 24800
rect 45787 24769 45799 24772
rect 45741 24763 45799 24769
rect 46293 24769 46305 24772
rect 46339 24800 46351 24803
rect 47026 24800 47032 24812
rect 46339 24772 47032 24800
rect 46339 24769 46351 24772
rect 46293 24763 46351 24769
rect 47026 24760 47032 24772
rect 47084 24760 47090 24812
rect 47762 24800 47768 24812
rect 47723 24772 47768 24800
rect 47762 24760 47768 24772
rect 47820 24760 47826 24812
rect 44358 24732 44364 24744
rect 39172 24704 40080 24732
rect 44319 24704 44364 24732
rect 39172 24692 39178 24704
rect 44358 24692 44364 24704
rect 44416 24692 44422 24744
rect 38010 24664 38016 24676
rect 36743 24636 38016 24664
rect 36633 24627 36691 24633
rect 38010 24624 38016 24636
rect 38068 24624 38074 24676
rect 45554 24664 45560 24676
rect 38948 24636 45560 24664
rect 24857 24599 24915 24605
rect 24857 24565 24869 24599
rect 24903 24596 24915 24599
rect 24946 24596 24952 24608
rect 24903 24568 24952 24596
rect 24903 24565 24915 24568
rect 24857 24559 24915 24565
rect 24946 24556 24952 24568
rect 25004 24556 25010 24608
rect 31113 24599 31171 24605
rect 31113 24565 31125 24599
rect 31159 24596 31171 24599
rect 31846 24596 31852 24608
rect 31159 24568 31852 24596
rect 31159 24565 31171 24568
rect 31113 24559 31171 24565
rect 31846 24556 31852 24568
rect 31904 24556 31910 24608
rect 34790 24556 34796 24608
rect 34848 24596 34854 24608
rect 35989 24599 36047 24605
rect 35989 24596 36001 24599
rect 34848 24568 36001 24596
rect 34848 24556 34854 24568
rect 35989 24565 36001 24568
rect 36035 24596 36047 24599
rect 36541 24599 36599 24605
rect 36541 24596 36553 24599
rect 36035 24568 36553 24596
rect 36035 24565 36047 24568
rect 35989 24559 36047 24565
rect 36541 24565 36553 24568
rect 36587 24565 36599 24599
rect 36541 24559 36599 24565
rect 37182 24556 37188 24608
rect 37240 24596 37246 24608
rect 38948 24596 38976 24636
rect 45554 24624 45560 24636
rect 45612 24624 45618 24676
rect 39390 24596 39396 24608
rect 37240 24568 38976 24596
rect 39351 24568 39396 24596
rect 37240 24556 37246 24568
rect 39390 24556 39396 24568
rect 39448 24556 39454 24608
rect 39853 24599 39911 24605
rect 39853 24565 39865 24599
rect 39899 24596 39911 24599
rect 40586 24596 40592 24608
rect 39899 24568 40592 24596
rect 39899 24565 39911 24568
rect 39853 24559 39911 24565
rect 40586 24556 40592 24568
rect 40644 24556 40650 24608
rect 44726 24596 44732 24608
rect 44687 24568 44732 24596
rect 44726 24556 44732 24568
rect 44784 24556 44790 24608
rect 45189 24599 45247 24605
rect 45189 24565 45201 24599
rect 45235 24596 45247 24599
rect 45462 24596 45468 24608
rect 45235 24568 45468 24596
rect 45235 24565 45247 24568
rect 45189 24559 45247 24565
rect 45462 24556 45468 24568
rect 45520 24556 45526 24608
rect 45830 24556 45836 24608
rect 45888 24596 45894 24608
rect 46385 24599 46443 24605
rect 46385 24596 46397 24599
rect 45888 24568 46397 24596
rect 45888 24556 45894 24568
rect 46385 24565 46397 24568
rect 46431 24565 46443 24599
rect 46385 24559 46443 24565
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 22097 24395 22155 24401
rect 22097 24361 22109 24395
rect 22143 24392 22155 24395
rect 22186 24392 22192 24404
rect 22143 24364 22192 24392
rect 22143 24361 22155 24364
rect 22097 24355 22155 24361
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 23290 24392 23296 24404
rect 23251 24364 23296 24392
rect 23290 24352 23296 24364
rect 23348 24352 23354 24404
rect 33686 24392 33692 24404
rect 24320 24364 33692 24392
rect 21910 24216 21916 24268
rect 21968 24256 21974 24268
rect 24320 24256 24348 24364
rect 33686 24352 33692 24364
rect 33744 24352 33750 24404
rect 38013 24395 38071 24401
rect 38013 24361 38025 24395
rect 38059 24392 38071 24395
rect 39025 24395 39083 24401
rect 39025 24392 39037 24395
rect 38059 24364 39037 24392
rect 38059 24361 38071 24364
rect 38013 24355 38071 24361
rect 39025 24361 39037 24364
rect 39071 24392 39083 24395
rect 39114 24392 39120 24404
rect 39071 24364 39120 24392
rect 39071 24361 39083 24364
rect 39025 24355 39083 24361
rect 39114 24352 39120 24364
rect 39172 24352 39178 24404
rect 39482 24352 39488 24404
rect 39540 24392 39546 24404
rect 39853 24395 39911 24401
rect 39853 24392 39865 24395
rect 39540 24364 39865 24392
rect 39540 24352 39546 24364
rect 39853 24361 39865 24364
rect 39899 24361 39911 24395
rect 39853 24355 39911 24361
rect 32122 24324 32128 24336
rect 21968 24228 24348 24256
rect 30392 24296 32128 24324
rect 21968 24216 21974 24228
rect 2038 24148 2044 24200
rect 2096 24188 2102 24200
rect 22020 24197 22048 24228
rect 2317 24191 2375 24197
rect 2317 24188 2329 24191
rect 2096 24160 2329 24188
rect 2096 24148 2102 24160
rect 2317 24157 2329 24160
rect 2363 24157 2375 24191
rect 2317 24151 2375 24157
rect 22005 24191 22063 24197
rect 22005 24157 22017 24191
rect 22051 24157 22063 24191
rect 22922 24188 22928 24200
rect 22883 24160 22928 24188
rect 22005 24151 22063 24157
rect 22922 24148 22928 24160
rect 22980 24148 22986 24200
rect 23385 24191 23443 24197
rect 23385 24157 23397 24191
rect 23431 24188 23443 24191
rect 23934 24188 23940 24200
rect 23431 24160 23940 24188
rect 23431 24157 23443 24160
rect 23385 24151 23443 24157
rect 23934 24148 23940 24160
rect 23992 24148 23998 24200
rect 24397 24191 24455 24197
rect 24397 24157 24409 24191
rect 24443 24188 24455 24191
rect 27617 24191 27675 24197
rect 24443 24160 24900 24188
rect 24443 24157 24455 24160
rect 24397 24151 24455 24157
rect 24872 24132 24900 24160
rect 27617 24157 27629 24191
rect 27663 24188 27675 24191
rect 28810 24188 28816 24200
rect 27663 24160 28816 24188
rect 27663 24157 27675 24160
rect 27617 24151 27675 24157
rect 28810 24148 28816 24160
rect 28868 24148 28874 24200
rect 30392 24197 30420 24296
rect 32122 24284 32128 24296
rect 32180 24284 32186 24336
rect 33134 24284 33140 24336
rect 33192 24324 33198 24336
rect 33962 24324 33968 24336
rect 33192 24296 33968 24324
rect 33192 24284 33198 24296
rect 33962 24284 33968 24296
rect 34020 24284 34026 24336
rect 40034 24324 40040 24336
rect 38212 24296 40040 24324
rect 30469 24259 30527 24265
rect 30469 24225 30481 24259
rect 30515 24256 30527 24259
rect 31110 24256 31116 24268
rect 30515 24228 31116 24256
rect 30515 24225 30527 24228
rect 30469 24219 30527 24225
rect 31110 24216 31116 24228
rect 31168 24256 31174 24268
rect 31168 24228 31616 24256
rect 31168 24216 31174 24228
rect 30377 24191 30435 24197
rect 30377 24157 30389 24191
rect 30423 24157 30435 24191
rect 31478 24188 31484 24200
rect 31439 24160 31484 24188
rect 30377 24151 30435 24157
rect 31478 24148 31484 24160
rect 31536 24148 31542 24200
rect 31588 24197 31616 24228
rect 32306 24216 32312 24268
rect 32364 24256 32370 24268
rect 34514 24256 34520 24268
rect 32364 24228 34520 24256
rect 32364 24216 32370 24228
rect 34514 24216 34520 24228
rect 34572 24256 34578 24268
rect 35434 24256 35440 24268
rect 34572 24228 35440 24256
rect 34572 24216 34578 24228
rect 35434 24216 35440 24228
rect 35492 24256 35498 24268
rect 35529 24259 35587 24265
rect 35529 24256 35541 24259
rect 35492 24228 35541 24256
rect 35492 24216 35498 24228
rect 35529 24225 35541 24228
rect 35575 24225 35587 24259
rect 35529 24219 35587 24225
rect 38010 24216 38016 24268
rect 38068 24256 38074 24268
rect 38212 24265 38240 24296
rect 40034 24284 40040 24296
rect 40092 24284 40098 24336
rect 46198 24324 46204 24336
rect 43088 24296 46204 24324
rect 38197 24259 38255 24265
rect 38197 24256 38209 24259
rect 38068 24228 38209 24256
rect 38068 24216 38074 24228
rect 38197 24225 38209 24228
rect 38243 24225 38255 24259
rect 38654 24256 38660 24268
rect 38197 24219 38255 24225
rect 38304 24228 38660 24256
rect 31573 24191 31631 24197
rect 31573 24157 31585 24191
rect 31619 24157 31631 24191
rect 31573 24151 31631 24157
rect 31662 24148 31668 24200
rect 31720 24188 31726 24200
rect 31757 24191 31815 24197
rect 31757 24188 31769 24191
rect 31720 24160 31769 24188
rect 31720 24148 31726 24160
rect 31757 24157 31769 24160
rect 31803 24157 31815 24191
rect 31757 24151 31815 24157
rect 31846 24148 31852 24200
rect 31904 24188 31910 24200
rect 32953 24191 33011 24197
rect 31904 24160 31949 24188
rect 31904 24148 31910 24160
rect 32953 24157 32965 24191
rect 32999 24157 33011 24191
rect 33134 24188 33140 24200
rect 33095 24160 33140 24188
rect 32953 24151 33011 24157
rect 22738 24080 22744 24132
rect 22796 24120 22802 24132
rect 23017 24123 23075 24129
rect 23017 24120 23029 24123
rect 22796 24092 23029 24120
rect 22796 24080 22802 24092
rect 23017 24089 23029 24092
rect 23063 24089 23075 24123
rect 24642 24123 24700 24129
rect 24642 24120 24654 24123
rect 23017 24083 23075 24089
rect 23400 24092 24654 24120
rect 23106 24052 23112 24064
rect 23067 24024 23112 24052
rect 23106 24012 23112 24024
rect 23164 24012 23170 24064
rect 23400 24061 23428 24092
rect 24642 24089 24654 24092
rect 24688 24089 24700 24123
rect 24642 24083 24700 24089
rect 24854 24080 24860 24132
rect 24912 24080 24918 24132
rect 27798 24080 27804 24132
rect 27856 24120 27862 24132
rect 28718 24120 28724 24132
rect 27856 24092 28724 24120
rect 27856 24080 27862 24092
rect 28718 24080 28724 24092
rect 28776 24080 28782 24132
rect 23385 24055 23443 24061
rect 23385 24021 23397 24055
rect 23431 24021 23443 24055
rect 23385 24015 23443 24021
rect 24762 24012 24768 24064
rect 24820 24052 24826 24064
rect 25777 24055 25835 24061
rect 25777 24052 25789 24055
rect 24820 24024 25789 24052
rect 24820 24012 24826 24024
rect 25777 24021 25789 24024
rect 25823 24021 25835 24055
rect 27982 24052 27988 24064
rect 27943 24024 27988 24052
rect 25777 24015 25835 24021
rect 27982 24012 27988 24024
rect 28040 24012 28046 24064
rect 30834 24012 30840 24064
rect 30892 24052 30898 24064
rect 31297 24055 31355 24061
rect 31297 24052 31309 24055
rect 30892 24024 31309 24052
rect 30892 24012 30898 24024
rect 31297 24021 31309 24024
rect 31343 24021 31355 24055
rect 32766 24052 32772 24064
rect 32727 24024 32772 24052
rect 31297 24015 31355 24021
rect 32766 24012 32772 24024
rect 32824 24012 32830 24064
rect 32968 24052 32996 24151
rect 33134 24148 33140 24160
rect 33192 24148 33198 24200
rect 33229 24191 33287 24197
rect 33229 24157 33241 24191
rect 33275 24188 33287 24191
rect 33594 24188 33600 24200
rect 33275 24160 33600 24188
rect 33275 24157 33287 24160
rect 33229 24151 33287 24157
rect 33594 24148 33600 24160
rect 33652 24188 33658 24200
rect 33873 24191 33931 24197
rect 33873 24188 33885 24191
rect 33652 24160 33885 24188
rect 33652 24148 33658 24160
rect 33873 24157 33885 24160
rect 33919 24157 33931 24191
rect 33873 24151 33931 24157
rect 33962 24148 33968 24200
rect 34020 24188 34026 24200
rect 34020 24160 34065 24188
rect 34020 24148 34026 24160
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 35802 24197 35808 24200
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 34848 24160 34897 24188
rect 34848 24148 34854 24160
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 35069 24191 35127 24197
rect 35069 24157 35081 24191
rect 35115 24157 35127 24191
rect 35796 24188 35808 24197
rect 35763 24160 35808 24188
rect 35069 24151 35127 24157
rect 35796 24151 35808 24160
rect 33318 24080 33324 24132
rect 33376 24120 33382 24132
rect 33689 24123 33747 24129
rect 33689 24120 33701 24123
rect 33376 24092 33701 24120
rect 33376 24080 33382 24092
rect 33689 24089 33701 24092
rect 33735 24089 33747 24123
rect 35084 24120 35112 24151
rect 35802 24148 35808 24151
rect 35860 24148 35866 24200
rect 37921 24191 37979 24197
rect 37921 24157 37933 24191
rect 37967 24188 37979 24191
rect 38304 24188 38332 24228
rect 38654 24216 38660 24228
rect 38712 24256 38718 24268
rect 39390 24256 39396 24268
rect 38712 24228 39396 24256
rect 38712 24216 38718 24228
rect 39390 24216 39396 24228
rect 39448 24216 39454 24268
rect 41414 24216 41420 24268
rect 41472 24256 41478 24268
rect 43088 24265 43116 24296
rect 46198 24284 46204 24296
rect 46256 24284 46262 24336
rect 43073 24259 43131 24265
rect 41472 24228 41517 24256
rect 41472 24216 41478 24228
rect 43073 24225 43085 24259
rect 43119 24225 43131 24259
rect 43073 24219 43131 24225
rect 43898 24216 43904 24268
rect 43956 24256 43962 24268
rect 46293 24259 46351 24265
rect 43956 24228 45324 24256
rect 43956 24216 43962 24228
rect 37967 24160 38332 24188
rect 37967 24157 37979 24160
rect 37921 24151 37979 24157
rect 38470 24148 38476 24200
rect 38528 24188 38534 24200
rect 38749 24191 38807 24197
rect 38749 24188 38761 24191
rect 38528 24160 38761 24188
rect 38528 24148 38534 24160
rect 38749 24157 38761 24160
rect 38795 24157 38807 24191
rect 38749 24151 38807 24157
rect 38841 24191 38899 24197
rect 38841 24157 38853 24191
rect 38887 24157 38899 24191
rect 38841 24151 38899 24157
rect 36262 24120 36268 24132
rect 33689 24083 33747 24089
rect 34808 24092 36268 24120
rect 34808 24064 34836 24092
rect 36262 24080 36268 24092
rect 36320 24080 36326 24132
rect 38194 24120 38200 24132
rect 38155 24092 38200 24120
rect 38194 24080 38200 24092
rect 38252 24080 38258 24132
rect 38378 24080 38384 24132
rect 38436 24120 38442 24132
rect 38856 24120 38884 24151
rect 39758 24148 39764 24200
rect 39816 24188 39822 24200
rect 39853 24191 39911 24197
rect 39853 24188 39865 24191
rect 39816 24160 39865 24188
rect 39816 24148 39822 24160
rect 39853 24157 39865 24160
rect 39899 24157 39911 24191
rect 39853 24151 39911 24157
rect 40037 24191 40095 24197
rect 40037 24157 40049 24191
rect 40083 24157 40095 24191
rect 41230 24188 41236 24200
rect 41191 24160 41236 24188
rect 40037 24151 40095 24157
rect 38436 24092 38884 24120
rect 38436 24080 38442 24092
rect 33787 24055 33845 24061
rect 33787 24052 33799 24055
rect 32968 24024 33799 24052
rect 33787 24021 33799 24024
rect 33833 24021 33845 24055
rect 33787 24015 33845 24021
rect 34790 24012 34796 24064
rect 34848 24012 34854 24064
rect 34977 24055 35035 24061
rect 34977 24021 34989 24055
rect 35023 24052 35035 24055
rect 35342 24052 35348 24064
rect 35023 24024 35348 24052
rect 35023 24021 35035 24024
rect 34977 24015 35035 24021
rect 35342 24012 35348 24024
rect 35400 24012 35406 24064
rect 36170 24012 36176 24064
rect 36228 24052 36234 24064
rect 36909 24055 36967 24061
rect 36909 24052 36921 24055
rect 36228 24024 36921 24052
rect 36228 24012 36234 24024
rect 36909 24021 36921 24024
rect 36955 24052 36967 24055
rect 37274 24052 37280 24064
rect 36955 24024 37280 24052
rect 36955 24021 36967 24024
rect 36909 24015 36967 24021
rect 37274 24012 37280 24024
rect 37332 24052 37338 24064
rect 37734 24052 37740 24064
rect 37332 24024 37740 24052
rect 37332 24012 37338 24024
rect 37734 24012 37740 24024
rect 37792 24012 37798 24064
rect 38838 24012 38844 24064
rect 38896 24052 38902 24064
rect 40052 24052 40080 24151
rect 41230 24148 41236 24160
rect 41288 24148 41294 24200
rect 43809 24191 43867 24197
rect 43809 24157 43821 24191
rect 43855 24157 43867 24191
rect 43990 24188 43996 24200
rect 43951 24160 43996 24188
rect 43809 24151 43867 24157
rect 43824 24120 43852 24151
rect 43990 24148 43996 24160
rect 44048 24148 44054 24200
rect 45189 24191 45247 24197
rect 45189 24157 45201 24191
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 44726 24120 44732 24132
rect 43824 24092 44732 24120
rect 44726 24080 44732 24092
rect 44784 24120 44790 24132
rect 45204 24120 45232 24151
rect 44784 24092 45232 24120
rect 45296 24120 45324 24228
rect 46293 24225 46305 24259
rect 46339 24256 46351 24259
rect 47762 24256 47768 24268
rect 46339 24228 47768 24256
rect 46339 24225 46351 24228
rect 46293 24219 46351 24225
rect 47762 24216 47768 24228
rect 47820 24216 47826 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 45462 24188 45468 24200
rect 45423 24160 45468 24188
rect 45462 24148 45468 24160
rect 45520 24148 45526 24200
rect 45373 24123 45431 24129
rect 45373 24120 45385 24123
rect 45296 24092 45385 24120
rect 44784 24080 44790 24092
rect 45373 24089 45385 24092
rect 45419 24089 45431 24123
rect 45373 24083 45431 24089
rect 46477 24123 46535 24129
rect 46477 24089 46489 24123
rect 46523 24120 46535 24123
rect 46934 24120 46940 24132
rect 46523 24092 46940 24120
rect 46523 24089 46535 24092
rect 46477 24083 46535 24089
rect 46934 24080 46940 24092
rect 46992 24080 46998 24132
rect 38896 24024 40080 24052
rect 38896 24012 38902 24024
rect 43806 24012 43812 24064
rect 43864 24052 43870 24064
rect 43901 24055 43959 24061
rect 43901 24052 43913 24055
rect 43864 24024 43913 24052
rect 43864 24012 43870 24024
rect 43901 24021 43913 24024
rect 43947 24021 43959 24055
rect 43901 24015 43959 24021
rect 45005 24055 45063 24061
rect 45005 24021 45017 24055
rect 45051 24052 45063 24055
rect 45094 24052 45100 24064
rect 45051 24024 45100 24052
rect 45051 24021 45063 24024
rect 45005 24015 45063 24021
rect 45094 24012 45100 24024
rect 45152 24012 45158 24064
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 22002 23808 22008 23860
rect 22060 23848 22066 23860
rect 24029 23851 24087 23857
rect 24029 23848 24041 23851
rect 22060 23820 24041 23848
rect 22060 23808 22066 23820
rect 24029 23817 24041 23820
rect 24075 23817 24087 23851
rect 27522 23848 27528 23860
rect 24029 23811 24087 23817
rect 25332 23820 27528 23848
rect 2038 23712 2044 23724
rect 1999 23684 2044 23712
rect 2038 23672 2044 23684
rect 2096 23672 2102 23724
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23681 24455 23715
rect 24397 23675 24455 23681
rect 24765 23715 24823 23721
rect 24765 23681 24777 23715
rect 24811 23712 24823 23715
rect 24946 23712 24952 23724
rect 24811 23684 24952 23712
rect 24811 23681 24823 23684
rect 24765 23675 24823 23681
rect 2222 23644 2228 23656
rect 2183 23616 2228 23644
rect 2222 23604 2228 23616
rect 2280 23604 2286 23656
rect 2774 23644 2780 23656
rect 2735 23616 2780 23644
rect 2774 23604 2780 23616
rect 2832 23604 2838 23656
rect 23934 23644 23940 23656
rect 23895 23616 23940 23644
rect 23934 23604 23940 23616
rect 23992 23604 23998 23656
rect 24302 23644 24308 23656
rect 24263 23616 24308 23644
rect 24302 23604 24308 23616
rect 24360 23604 24366 23656
rect 24412 23576 24440 23675
rect 24946 23672 24952 23684
rect 25004 23672 25010 23724
rect 24578 23604 24584 23656
rect 24636 23644 24642 23656
rect 24673 23647 24731 23653
rect 24673 23644 24685 23647
rect 24636 23616 24685 23644
rect 24636 23604 24642 23616
rect 24673 23613 24685 23616
rect 24719 23613 24731 23647
rect 25332 23644 25360 23820
rect 27522 23808 27528 23820
rect 27580 23808 27586 23860
rect 30374 23808 30380 23860
rect 30432 23848 30438 23860
rect 30432 23820 31432 23848
rect 30432 23808 30438 23820
rect 27709 23783 27767 23789
rect 27709 23780 27721 23783
rect 25424 23752 27721 23780
rect 25424 23721 25452 23752
rect 27709 23749 27721 23752
rect 27755 23749 27767 23783
rect 27709 23743 27767 23749
rect 28629 23783 28687 23789
rect 28629 23749 28641 23783
rect 28675 23780 28687 23783
rect 31202 23780 31208 23792
rect 28675 23752 31208 23780
rect 28675 23749 28687 23752
rect 28629 23743 28687 23749
rect 31202 23740 31208 23752
rect 31260 23740 31266 23792
rect 25409 23715 25467 23721
rect 25409 23681 25421 23715
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 25502 23715 25560 23721
rect 25502 23681 25514 23715
rect 25548 23681 25560 23715
rect 25682 23712 25688 23724
rect 25643 23684 25688 23712
rect 25502 23675 25560 23681
rect 25516 23644 25544 23675
rect 25682 23672 25688 23684
rect 25740 23672 25746 23724
rect 25774 23672 25780 23724
rect 25832 23712 25838 23724
rect 25958 23721 25964 23724
rect 25913 23715 25964 23721
rect 25832 23684 25874 23712
rect 25832 23672 25838 23684
rect 25913 23681 25925 23715
rect 25959 23681 25964 23715
rect 25913 23675 25964 23681
rect 25958 23672 25964 23675
rect 26016 23672 26022 23724
rect 26970 23712 26976 23724
rect 26931 23684 26976 23712
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 27154 23672 27160 23724
rect 27212 23714 27218 23724
rect 27212 23686 27255 23714
rect 27212 23672 27218 23686
rect 27522 23672 27528 23724
rect 27580 23712 27586 23724
rect 30834 23712 30840 23724
rect 27580 23684 27625 23712
rect 30795 23684 30840 23712
rect 27580 23672 27586 23684
rect 30834 23672 30840 23684
rect 30892 23672 30898 23724
rect 31018 23712 31024 23724
rect 30979 23684 31024 23712
rect 31018 23672 31024 23684
rect 31076 23672 31082 23724
rect 31110 23672 31116 23724
rect 31168 23712 31174 23724
rect 31404 23721 31432 23820
rect 33594 23808 33600 23860
rect 33652 23848 33658 23860
rect 33873 23851 33931 23857
rect 33873 23848 33885 23851
rect 33652 23820 33885 23848
rect 33652 23808 33658 23820
rect 33873 23817 33885 23820
rect 33919 23817 33931 23851
rect 33873 23811 33931 23817
rect 35986 23808 35992 23860
rect 36044 23848 36050 23860
rect 36541 23851 36599 23857
rect 36541 23848 36553 23851
rect 36044 23820 36553 23848
rect 36044 23808 36050 23820
rect 36541 23817 36553 23820
rect 36587 23817 36599 23851
rect 36541 23811 36599 23817
rect 38378 23808 38384 23860
rect 38436 23848 38442 23860
rect 38673 23851 38731 23857
rect 38673 23848 38685 23851
rect 38436 23820 38685 23848
rect 38436 23808 38442 23820
rect 38673 23817 38685 23820
rect 38719 23817 38731 23851
rect 38838 23848 38844 23860
rect 38799 23820 38844 23848
rect 38673 23811 38731 23817
rect 38838 23808 38844 23820
rect 38896 23808 38902 23860
rect 39574 23848 39580 23860
rect 39535 23820 39580 23848
rect 39574 23808 39580 23820
rect 39632 23808 39638 23860
rect 43165 23851 43223 23857
rect 43165 23817 43177 23851
rect 43211 23848 43223 23851
rect 43990 23848 43996 23860
rect 43211 23820 43996 23848
rect 43211 23817 43223 23820
rect 43165 23811 43223 23817
rect 43990 23808 43996 23820
rect 44048 23808 44054 23860
rect 46934 23848 46940 23860
rect 46895 23820 46940 23848
rect 46934 23808 46940 23820
rect 46992 23808 46998 23860
rect 32766 23789 32772 23792
rect 32760 23780 32772 23789
rect 32727 23752 32772 23780
rect 32760 23743 32772 23752
rect 32766 23740 32772 23743
rect 32824 23740 32830 23792
rect 36170 23740 36176 23792
rect 36228 23780 36234 23792
rect 36389 23783 36447 23789
rect 36389 23780 36401 23783
rect 36228 23752 36273 23780
rect 36228 23740 36234 23752
rect 36372 23749 36401 23780
rect 36435 23780 36447 23783
rect 38473 23783 38531 23789
rect 36435 23752 37320 23780
rect 36435 23749 36447 23752
rect 36372 23743 36447 23749
rect 31389 23715 31447 23721
rect 31168 23684 31213 23712
rect 31168 23672 31174 23684
rect 31389 23681 31401 23715
rect 31435 23681 31447 23715
rect 31389 23675 31447 23681
rect 32306 23672 32312 23724
rect 32364 23712 32370 23724
rect 32493 23715 32551 23721
rect 32493 23712 32505 23715
rect 32364 23684 32505 23712
rect 32364 23672 32370 23684
rect 32493 23681 32505 23684
rect 32539 23681 32551 23715
rect 32493 23675 32551 23681
rect 34333 23715 34391 23721
rect 34333 23681 34345 23715
rect 34379 23712 34391 23715
rect 34422 23712 34428 23724
rect 34379 23684 34428 23712
rect 34379 23681 34391 23684
rect 34333 23675 34391 23681
rect 34422 23672 34428 23684
rect 34480 23672 34486 23724
rect 34606 23721 34612 23724
rect 34600 23675 34612 23721
rect 34664 23712 34670 23724
rect 34664 23684 34700 23712
rect 34606 23672 34612 23675
rect 34664 23672 34670 23684
rect 35710 23672 35716 23724
rect 35768 23712 35774 23724
rect 36372 23712 36400 23743
rect 35768 23684 36400 23712
rect 37292 23712 37320 23752
rect 38473 23749 38485 23783
rect 38519 23780 38531 23783
rect 38562 23780 38568 23792
rect 38519 23752 38568 23780
rect 38519 23749 38531 23752
rect 38473 23743 38531 23749
rect 38562 23740 38568 23752
rect 38620 23740 38626 23792
rect 38856 23712 38884 23808
rect 42426 23780 42432 23792
rect 40512 23752 42432 23780
rect 37292 23684 38884 23712
rect 39301 23715 39359 23721
rect 35768 23672 35774 23684
rect 39301 23681 39313 23715
rect 39347 23712 39359 23715
rect 39347 23684 39528 23712
rect 39347 23681 39359 23684
rect 39301 23675 39359 23681
rect 27243 23647 27301 23653
rect 27243 23644 27255 23647
rect 25332 23616 25544 23644
rect 27080 23616 27255 23644
rect 24673 23607 24731 23613
rect 26053 23579 26111 23585
rect 26053 23576 26065 23579
rect 24412 23548 26065 23576
rect 26053 23545 26065 23548
rect 26099 23545 26111 23579
rect 26053 23539 26111 23545
rect 26786 23536 26792 23588
rect 26844 23576 26850 23588
rect 27080 23576 27108 23616
rect 27243 23613 27255 23616
rect 27289 23613 27301 23647
rect 27243 23607 27301 23613
rect 27341 23647 27399 23653
rect 27341 23613 27353 23647
rect 27387 23644 27399 23647
rect 27387 23616 27476 23644
rect 27387 23613 27399 23616
rect 27341 23607 27399 23613
rect 26844 23548 27108 23576
rect 26844 23536 26850 23548
rect 25682 23468 25688 23520
rect 25740 23508 25746 23520
rect 26418 23508 26424 23520
rect 25740 23480 26424 23508
rect 25740 23468 25746 23480
rect 26418 23468 26424 23480
rect 26476 23508 26482 23520
rect 27448 23508 27476 23616
rect 30742 23604 30748 23656
rect 30800 23644 30806 23656
rect 31205 23647 31263 23653
rect 31205 23644 31217 23647
rect 30800 23616 31217 23644
rect 30800 23604 30806 23616
rect 31205 23613 31217 23616
rect 31251 23613 31263 23647
rect 31205 23607 31263 23613
rect 38378 23536 38384 23588
rect 38436 23576 38442 23588
rect 39393 23579 39451 23585
rect 39393 23576 39405 23579
rect 38436 23548 39405 23576
rect 38436 23536 38442 23548
rect 39393 23545 39405 23548
rect 39439 23545 39451 23579
rect 39393 23539 39451 23545
rect 39500 23576 39528 23684
rect 39850 23672 39856 23724
rect 39908 23712 39914 23724
rect 40512 23721 40540 23752
rect 42426 23740 42432 23752
rect 42484 23740 42490 23792
rect 43272 23752 44588 23780
rect 43272 23724 43300 23752
rect 40497 23715 40555 23721
rect 40497 23712 40509 23715
rect 39908 23684 40509 23712
rect 39908 23672 39914 23684
rect 40497 23681 40509 23684
rect 40543 23681 40555 23715
rect 40497 23675 40555 23681
rect 40586 23672 40592 23724
rect 40644 23712 40650 23724
rect 40753 23715 40811 23721
rect 40753 23712 40765 23715
rect 40644 23684 40765 23712
rect 40644 23672 40650 23684
rect 40753 23681 40765 23684
rect 40799 23681 40811 23715
rect 40753 23675 40811 23681
rect 43073 23715 43131 23721
rect 43073 23681 43085 23715
rect 43119 23712 43131 23715
rect 43162 23712 43168 23724
rect 43119 23684 43168 23712
rect 43119 23681 43131 23684
rect 43073 23675 43131 23681
rect 43162 23672 43168 23684
rect 43220 23672 43226 23724
rect 43254 23672 43260 23724
rect 43312 23712 43318 23724
rect 43898 23712 43904 23724
rect 43312 23684 43357 23712
rect 43640 23684 43904 23712
rect 43312 23672 43318 23684
rect 39577 23647 39635 23653
rect 39577 23613 39589 23647
rect 39623 23644 39635 23647
rect 40034 23644 40040 23656
rect 39623 23616 40040 23644
rect 39623 23613 39635 23616
rect 39577 23607 39635 23613
rect 40034 23604 40040 23616
rect 40092 23604 40098 23656
rect 42794 23604 42800 23656
rect 42852 23644 42858 23656
rect 43640 23644 43668 23684
rect 43898 23672 43904 23684
rect 43956 23672 43962 23724
rect 44560 23712 44588 23752
rect 45830 23712 45836 23724
rect 44560 23684 45836 23712
rect 45830 23672 45836 23684
rect 45888 23721 45894 23724
rect 45888 23715 45937 23721
rect 45888 23681 45891 23715
rect 45925 23681 45937 23715
rect 46014 23712 46020 23724
rect 45975 23684 46020 23712
rect 45888 23675 45937 23681
rect 45888 23672 45894 23675
rect 46014 23672 46020 23684
rect 46072 23672 46078 23724
rect 46106 23672 46112 23724
rect 46164 23712 46170 23724
rect 46164 23684 46209 23712
rect 46164 23672 46170 23684
rect 46290 23672 46296 23724
rect 46348 23712 46354 23724
rect 46845 23715 46903 23721
rect 46348 23684 46393 23712
rect 46348 23672 46354 23684
rect 46845 23681 46857 23715
rect 46891 23712 46903 23715
rect 47210 23712 47216 23724
rect 46891 23684 47216 23712
rect 46891 23681 46903 23684
rect 46845 23675 46903 23681
rect 47210 23672 47216 23684
rect 47268 23672 47274 23724
rect 47762 23712 47768 23724
rect 47723 23684 47768 23712
rect 47762 23672 47768 23684
rect 47820 23672 47826 23724
rect 43806 23644 43812 23656
rect 42852 23616 43668 23644
rect 43767 23616 43812 23644
rect 42852 23604 42858 23616
rect 43806 23604 43812 23616
rect 43864 23604 43870 23656
rect 44269 23579 44327 23585
rect 39500 23548 39896 23576
rect 26476 23480 27476 23508
rect 26476 23468 26482 23480
rect 29546 23468 29552 23520
rect 29604 23508 29610 23520
rect 29917 23511 29975 23517
rect 29917 23508 29929 23511
rect 29604 23480 29929 23508
rect 29604 23468 29610 23480
rect 29917 23477 29929 23480
rect 29963 23477 29975 23511
rect 29917 23471 29975 23477
rect 30006 23468 30012 23520
rect 30064 23508 30070 23520
rect 31573 23511 31631 23517
rect 31573 23508 31585 23511
rect 30064 23480 31585 23508
rect 30064 23468 30070 23480
rect 31573 23477 31585 23480
rect 31619 23477 31631 23511
rect 31573 23471 31631 23477
rect 35526 23468 35532 23520
rect 35584 23508 35590 23520
rect 35713 23511 35771 23517
rect 35713 23508 35725 23511
rect 35584 23480 35725 23508
rect 35584 23468 35590 23480
rect 35713 23477 35725 23480
rect 35759 23508 35771 23511
rect 36357 23511 36415 23517
rect 36357 23508 36369 23511
rect 35759 23480 36369 23508
rect 35759 23477 35771 23480
rect 35713 23471 35771 23477
rect 36357 23477 36369 23480
rect 36403 23508 36415 23511
rect 36630 23508 36636 23520
rect 36403 23480 36636 23508
rect 36403 23477 36415 23480
rect 36357 23471 36415 23477
rect 36630 23468 36636 23480
rect 36688 23468 36694 23520
rect 38470 23468 38476 23520
rect 38528 23508 38534 23520
rect 38657 23511 38715 23517
rect 38657 23508 38669 23511
rect 38528 23480 38669 23508
rect 38528 23468 38534 23480
rect 38657 23477 38669 23480
rect 38703 23508 38715 23511
rect 39500 23508 39528 23548
rect 39868 23520 39896 23548
rect 44269 23545 44281 23579
rect 44315 23576 44327 23579
rect 45002 23576 45008 23588
rect 44315 23548 45008 23576
rect 44315 23545 44327 23548
rect 44269 23539 44327 23545
rect 45002 23536 45008 23548
rect 45060 23536 45066 23588
rect 38703 23480 39528 23508
rect 38703 23477 38715 23480
rect 38657 23471 38715 23477
rect 39850 23468 39856 23520
rect 39908 23508 39914 23520
rect 41877 23511 41935 23517
rect 41877 23508 41889 23511
rect 39908 23480 41889 23508
rect 39908 23468 39914 23480
rect 41877 23477 41889 23480
rect 41923 23477 41935 23511
rect 41877 23471 41935 23477
rect 45649 23511 45707 23517
rect 45649 23477 45661 23511
rect 45695 23508 45707 23511
rect 46934 23508 46940 23520
rect 45695 23480 46940 23508
rect 45695 23477 45707 23480
rect 45649 23471 45707 23477
rect 46934 23468 46940 23480
rect 46992 23468 46998 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 2222 23264 2228 23316
rect 2280 23304 2286 23316
rect 2409 23307 2467 23313
rect 2409 23304 2421 23307
rect 2280 23276 2421 23304
rect 2280 23264 2286 23276
rect 2409 23273 2421 23276
rect 2455 23273 2467 23307
rect 2409 23267 2467 23273
rect 24302 23264 24308 23316
rect 24360 23304 24366 23316
rect 24397 23307 24455 23313
rect 24397 23304 24409 23307
rect 24360 23276 24409 23304
rect 24360 23264 24366 23276
rect 24397 23273 24409 23276
rect 24443 23273 24455 23307
rect 24397 23267 24455 23273
rect 26970 23264 26976 23316
rect 27028 23304 27034 23316
rect 27801 23307 27859 23313
rect 27801 23304 27813 23307
rect 27028 23276 27813 23304
rect 27028 23264 27034 23276
rect 27801 23273 27813 23276
rect 27847 23273 27859 23307
rect 27801 23267 27859 23273
rect 32306 23264 32312 23316
rect 32364 23304 32370 23316
rect 32493 23307 32551 23313
rect 32493 23304 32505 23307
rect 32364 23276 32505 23304
rect 32364 23264 32370 23276
rect 32493 23273 32505 23276
rect 32539 23273 32551 23307
rect 32493 23267 32551 23273
rect 34606 23264 34612 23316
rect 34664 23304 34670 23316
rect 35069 23307 35127 23313
rect 35069 23304 35081 23307
rect 34664 23276 35081 23304
rect 34664 23264 34670 23276
rect 35069 23273 35081 23276
rect 35115 23273 35127 23307
rect 35069 23267 35127 23273
rect 35437 23307 35495 23313
rect 35437 23273 35449 23307
rect 35483 23304 35495 23307
rect 35710 23304 35716 23316
rect 35483 23276 35716 23304
rect 35483 23273 35495 23276
rect 35437 23267 35495 23273
rect 35710 23264 35716 23276
rect 35768 23264 35774 23316
rect 36906 23304 36912 23316
rect 36648 23276 36912 23304
rect 24578 23196 24584 23248
rect 24636 23236 24642 23248
rect 24857 23239 24915 23245
rect 24857 23236 24869 23239
rect 24636 23208 24869 23236
rect 24636 23196 24642 23208
rect 24857 23205 24869 23208
rect 24903 23205 24915 23239
rect 28997 23239 29055 23245
rect 28997 23236 29009 23239
rect 24857 23199 24915 23205
rect 27264 23208 29009 23236
rect 22094 23128 22100 23180
rect 22152 23168 22158 23180
rect 25774 23168 25780 23180
rect 22152 23140 25780 23168
rect 22152 23128 22158 23140
rect 2222 23060 2228 23112
rect 2280 23100 2286 23112
rect 2317 23103 2375 23109
rect 2317 23100 2329 23103
rect 2280 23072 2329 23100
rect 2280 23060 2286 23072
rect 2317 23069 2329 23072
rect 2363 23100 2375 23103
rect 16942 23100 16948 23112
rect 2363 23072 16948 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 16942 23060 16948 23072
rect 17000 23060 17006 23112
rect 24688 23109 24716 23140
rect 25774 23128 25780 23140
rect 25832 23128 25838 23180
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 24673 23103 24731 23109
rect 24673 23069 24685 23103
rect 24719 23069 24731 23103
rect 24946 23100 24952 23112
rect 24907 23072 24952 23100
rect 24673 23063 24731 23069
rect 24596 23032 24624 23063
rect 24946 23060 24952 23072
rect 25004 23060 25010 23112
rect 27264 23109 27292 23208
rect 28997 23205 29009 23208
rect 29043 23205 29055 23239
rect 30466 23236 30472 23248
rect 30427 23208 30472 23236
rect 28997 23199 29055 23205
rect 30466 23196 30472 23208
rect 30524 23196 30530 23248
rect 30650 23196 30656 23248
rect 30708 23236 30714 23248
rect 36648 23236 36676 23276
rect 36906 23264 36912 23276
rect 36964 23304 36970 23316
rect 41138 23304 41144 23316
rect 36964 23276 41144 23304
rect 36964 23264 36970 23276
rect 41138 23264 41144 23276
rect 41196 23264 41202 23316
rect 41230 23264 41236 23316
rect 41288 23304 41294 23316
rect 41325 23307 41383 23313
rect 41325 23304 41337 23307
rect 41288 23276 41337 23304
rect 41288 23264 41294 23276
rect 41325 23273 41337 23276
rect 41371 23273 41383 23307
rect 41325 23267 41383 23273
rect 45097 23307 45155 23313
rect 45097 23273 45109 23307
rect 45143 23304 45155 23307
rect 46106 23304 46112 23316
rect 45143 23276 46112 23304
rect 45143 23273 45155 23276
rect 45097 23267 45155 23273
rect 46106 23264 46112 23276
rect 46164 23264 46170 23316
rect 47026 23264 47032 23316
rect 47084 23304 47090 23316
rect 48041 23307 48099 23313
rect 48041 23304 48053 23307
rect 47084 23276 48053 23304
rect 47084 23264 47090 23276
rect 48041 23273 48053 23276
rect 48087 23273 48099 23307
rect 48041 23267 48099 23273
rect 30708 23208 36676 23236
rect 30708 23196 30714 23208
rect 39758 23196 39764 23248
rect 39816 23236 39822 23248
rect 39816 23208 41184 23236
rect 39816 23196 39822 23208
rect 27982 23168 27988 23180
rect 27448 23140 27988 23168
rect 27448 23109 27476 23140
rect 27982 23128 27988 23140
rect 28040 23128 28046 23180
rect 30006 23168 30012 23180
rect 28368 23140 30012 23168
rect 28368 23109 28396 23140
rect 30006 23128 30012 23140
rect 30064 23128 30070 23180
rect 39022 23168 39028 23180
rect 31726 23140 39028 23168
rect 27249 23103 27307 23109
rect 27249 23069 27261 23103
rect 27295 23069 27307 23103
rect 27249 23063 27307 23069
rect 27433 23103 27491 23109
rect 27433 23069 27445 23103
rect 27479 23069 27491 23103
rect 27433 23063 27491 23069
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23069 27675 23103
rect 27617 23063 27675 23069
rect 28353 23103 28411 23109
rect 28353 23069 28365 23103
rect 28399 23069 28411 23103
rect 28353 23063 28411 23069
rect 28501 23103 28559 23109
rect 28501 23069 28513 23103
rect 28547 23100 28559 23103
rect 28718 23100 28724 23112
rect 28547 23069 28580 23100
rect 28679 23072 28724 23100
rect 28501 23063 28580 23069
rect 25774 23032 25780 23044
rect 24596 23004 25780 23032
rect 25774 22992 25780 23004
rect 25832 22992 25838 23044
rect 26786 22992 26792 23044
rect 26844 23032 26850 23044
rect 27525 23035 27583 23041
rect 27525 23032 27537 23035
rect 26844 23004 27537 23032
rect 26844 22992 26850 23004
rect 27525 23001 27537 23004
rect 27571 23001 27583 23035
rect 27525 22995 27583 23001
rect 27154 22924 27160 22976
rect 27212 22964 27218 22976
rect 27430 22964 27436 22976
rect 27212 22936 27436 22964
rect 27212 22924 27218 22936
rect 27430 22924 27436 22936
rect 27488 22964 27494 22976
rect 27632 22964 27660 23063
rect 27488 22936 27660 22964
rect 28552 22964 28580 23063
rect 28718 23060 28724 23072
rect 28776 23060 28782 23112
rect 28810 23060 28816 23112
rect 28868 23109 28874 23112
rect 28868 23100 28876 23109
rect 30558 23100 30564 23112
rect 28868 23072 28913 23100
rect 30208 23072 30564 23100
rect 28868 23063 28876 23072
rect 28868 23060 28874 23063
rect 28629 23035 28687 23041
rect 28629 23001 28641 23035
rect 28675 23032 28687 23035
rect 30208 23032 30236 23072
rect 30558 23060 30564 23072
rect 30616 23060 30622 23112
rect 30745 23103 30803 23109
rect 30745 23069 30757 23103
rect 30791 23100 30803 23103
rect 31018 23100 31024 23112
rect 30791 23072 31024 23100
rect 30791 23069 30803 23072
rect 30745 23063 30803 23069
rect 31018 23060 31024 23072
rect 31076 23060 31082 23112
rect 31202 23100 31208 23112
rect 31163 23072 31208 23100
rect 31202 23060 31208 23072
rect 31260 23100 31266 23112
rect 31726 23100 31754 23140
rect 39022 23128 39028 23140
rect 39080 23128 39086 23180
rect 31260 23072 31754 23100
rect 35253 23103 35311 23109
rect 31260 23060 31266 23072
rect 35253 23069 35265 23103
rect 35299 23100 35311 23103
rect 35342 23100 35348 23112
rect 35299 23072 35348 23100
rect 35299 23069 35311 23072
rect 35253 23063 35311 23069
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 35526 23060 35532 23112
rect 35584 23100 35590 23112
rect 36265 23103 36323 23109
rect 35584 23072 35629 23100
rect 35584 23060 35590 23072
rect 36265 23069 36277 23103
rect 36311 23100 36323 23103
rect 36446 23100 36452 23112
rect 36311 23072 36452 23100
rect 36311 23069 36323 23072
rect 36265 23063 36323 23069
rect 36446 23060 36452 23072
rect 36504 23060 36510 23112
rect 37734 23100 37740 23112
rect 37695 23072 37740 23100
rect 37734 23060 37740 23072
rect 37792 23060 37798 23112
rect 39850 23100 39856 23112
rect 39811 23072 39856 23100
rect 39850 23060 39856 23072
rect 39908 23060 39914 23112
rect 39942 23060 39948 23112
rect 40000 23060 40006 23112
rect 40586 23100 40592 23112
rect 40547 23072 40592 23100
rect 40586 23060 40592 23072
rect 40644 23060 40650 23112
rect 40770 23100 40776 23112
rect 40731 23072 40776 23100
rect 40770 23060 40776 23072
rect 40828 23060 40834 23112
rect 41156 23109 41184 23208
rect 40865 23103 40923 23109
rect 40865 23069 40877 23103
rect 40911 23069 40923 23103
rect 40865 23063 40923 23069
rect 40957 23103 41015 23109
rect 40957 23069 40969 23103
rect 41003 23069 41015 23103
rect 40957 23063 41015 23069
rect 41141 23103 41199 23109
rect 41141 23069 41153 23103
rect 41187 23069 41199 23103
rect 45002 23100 45008 23112
rect 44963 23072 45008 23100
rect 41141 23063 41199 23069
rect 28675 23004 30236 23032
rect 28675 23001 28687 23004
rect 28629 22995 28687 23001
rect 30282 22992 30288 23044
rect 30340 23032 30346 23044
rect 30469 23035 30527 23041
rect 30469 23032 30481 23035
rect 30340 23004 30481 23032
rect 30340 22992 30346 23004
rect 30469 23001 30481 23004
rect 30515 23032 30527 23035
rect 39960 23032 39988 23060
rect 30515 23004 31754 23032
rect 30515 23001 30527 23004
rect 30469 22995 30527 23001
rect 30374 22964 30380 22976
rect 28552 22936 30380 22964
rect 27488 22924 27494 22936
rect 30374 22924 30380 22936
rect 30432 22924 30438 22976
rect 30558 22924 30564 22976
rect 30616 22964 30622 22976
rect 30653 22967 30711 22973
rect 30653 22964 30665 22967
rect 30616 22936 30665 22964
rect 30616 22924 30622 22936
rect 30653 22933 30665 22936
rect 30699 22933 30711 22967
rect 31726 22964 31754 23004
rect 39500 23004 39988 23032
rect 39500 22976 39528 23004
rect 40034 22992 40040 23044
rect 40092 23032 40098 23044
rect 40880 23032 40908 23063
rect 40092 23004 40908 23032
rect 40092 22992 40098 23004
rect 35894 22964 35900 22976
rect 31726 22936 35900 22964
rect 30653 22927 30711 22933
rect 35894 22924 35900 22936
rect 35952 22964 35958 22976
rect 36357 22967 36415 22973
rect 36357 22964 36369 22967
rect 35952 22936 36369 22964
rect 35952 22924 35958 22936
rect 36357 22933 36369 22936
rect 36403 22933 36415 22967
rect 36357 22927 36415 22933
rect 37829 22967 37887 22973
rect 37829 22933 37841 22967
rect 37875 22964 37887 22967
rect 39482 22964 39488 22976
rect 37875 22936 39488 22964
rect 37875 22933 37887 22936
rect 37829 22927 37887 22933
rect 39482 22924 39488 22936
rect 39540 22924 39546 22976
rect 39574 22924 39580 22976
rect 39632 22964 39638 22976
rect 39945 22967 40003 22973
rect 39945 22964 39957 22967
rect 39632 22936 39957 22964
rect 39632 22924 39638 22936
rect 39945 22933 39957 22936
rect 39991 22933 40003 22967
rect 39945 22927 40003 22933
rect 40126 22924 40132 22976
rect 40184 22964 40190 22976
rect 40972 22964 41000 23063
rect 45002 23060 45008 23072
rect 45060 23060 45066 23112
rect 45189 23103 45247 23109
rect 45189 23069 45201 23103
rect 45235 23100 45247 23103
rect 45278 23100 45284 23112
rect 45235 23072 45284 23100
rect 45235 23069 45247 23072
rect 45189 23063 45247 23069
rect 45278 23060 45284 23072
rect 45336 23060 45342 23112
rect 45646 23060 45652 23112
rect 45704 23100 45710 23112
rect 46658 23100 46664 23112
rect 45704 23072 46664 23100
rect 45704 23060 45710 23072
rect 46658 23060 46664 23072
rect 46716 23060 46722 23112
rect 46934 23109 46940 23112
rect 46928 23100 46940 23109
rect 46895 23072 46940 23100
rect 46928 23063 46940 23072
rect 46934 23060 46940 23063
rect 46992 23060 46998 23112
rect 40184 22936 41000 22964
rect 40184 22924 40190 22936
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 17862 22720 17868 22772
rect 17920 22760 17926 22772
rect 30650 22760 30656 22772
rect 17920 22732 30656 22760
rect 17920 22720 17926 22732
rect 30650 22720 30656 22732
rect 30708 22720 30714 22772
rect 30929 22763 30987 22769
rect 30929 22729 30941 22763
rect 30975 22760 30987 22763
rect 31018 22760 31024 22772
rect 30975 22732 31024 22760
rect 30975 22729 30987 22732
rect 30929 22723 30987 22729
rect 31018 22720 31024 22732
rect 31076 22760 31082 22772
rect 31478 22760 31484 22772
rect 31076 22732 31484 22760
rect 31076 22720 31082 22732
rect 31478 22720 31484 22732
rect 31536 22720 31542 22772
rect 33134 22760 33140 22772
rect 32416 22732 33140 22760
rect 23934 22652 23940 22704
rect 23992 22692 23998 22704
rect 24397 22695 24455 22701
rect 24397 22692 24409 22695
rect 23992 22664 24409 22692
rect 23992 22652 23998 22664
rect 24397 22661 24409 22664
rect 24443 22692 24455 22695
rect 30282 22692 30288 22704
rect 24443 22664 30288 22692
rect 24443 22661 24455 22664
rect 24397 22655 24455 22661
rect 30282 22652 30288 22664
rect 30340 22652 30346 22704
rect 24578 22624 24584 22636
rect 24539 22596 24584 22624
rect 24578 22584 24584 22596
rect 24636 22584 24642 22636
rect 24670 22584 24676 22636
rect 24728 22624 24734 22636
rect 29546 22624 29552 22636
rect 24728 22596 24773 22624
rect 29507 22596 29552 22624
rect 24728 22584 24734 22596
rect 29546 22584 29552 22596
rect 29604 22584 29610 22636
rect 29822 22633 29828 22636
rect 29816 22587 29828 22633
rect 29880 22624 29886 22636
rect 31573 22627 31631 22633
rect 29880 22596 29916 22624
rect 29822 22584 29828 22587
rect 29880 22584 29886 22596
rect 31573 22593 31585 22627
rect 31619 22624 31631 22627
rect 31662 22624 31668 22636
rect 31619 22596 31668 22624
rect 31619 22593 31631 22596
rect 31573 22587 31631 22593
rect 31662 22584 31668 22596
rect 31720 22584 31726 22636
rect 32416 22633 32444 22732
rect 33134 22720 33140 22732
rect 33192 22720 33198 22772
rect 33410 22720 33416 22772
rect 33468 22760 33474 22772
rect 34425 22763 34483 22769
rect 34425 22760 34437 22763
rect 33468 22732 34437 22760
rect 33468 22720 33474 22732
rect 34425 22729 34437 22732
rect 34471 22729 34483 22763
rect 34425 22723 34483 22729
rect 38013 22763 38071 22769
rect 38013 22729 38025 22763
rect 38059 22760 38071 22763
rect 39853 22763 39911 22769
rect 38059 22732 39712 22760
rect 38059 22729 38071 22732
rect 38013 22723 38071 22729
rect 32493 22695 32551 22701
rect 32493 22661 32505 22695
rect 32539 22692 32551 22695
rect 33290 22695 33348 22701
rect 33290 22692 33302 22695
rect 32539 22664 33302 22692
rect 32539 22661 32551 22664
rect 32493 22655 32551 22661
rect 33290 22661 33302 22664
rect 33336 22661 33348 22695
rect 35894 22692 35900 22704
rect 35855 22664 35900 22692
rect 33290 22655 33348 22661
rect 35894 22652 35900 22664
rect 35952 22652 35958 22704
rect 36081 22695 36139 22701
rect 36081 22661 36093 22695
rect 36127 22692 36139 22695
rect 37182 22692 37188 22704
rect 36127 22664 37188 22692
rect 36127 22661 36139 22664
rect 36081 22655 36139 22661
rect 37182 22652 37188 22664
rect 37240 22692 37246 22704
rect 39482 22692 39488 22704
rect 37240 22664 37964 22692
rect 39443 22664 39488 22692
rect 37240 22652 37246 22664
rect 32401 22627 32459 22633
rect 32401 22593 32413 22627
rect 32447 22593 32459 22627
rect 32582 22624 32588 22636
rect 32543 22596 32588 22624
rect 32401 22587 32459 22593
rect 32582 22584 32588 22596
rect 32640 22584 32646 22636
rect 35986 22584 35992 22636
rect 36044 22624 36050 22636
rect 36173 22627 36231 22633
rect 36173 22624 36185 22627
rect 36044 22596 36185 22624
rect 36044 22584 36050 22596
rect 36173 22593 36185 22596
rect 36219 22624 36231 22627
rect 36538 22624 36544 22636
rect 36219 22596 36544 22624
rect 36219 22593 36231 22596
rect 36173 22587 36231 22593
rect 36538 22584 36544 22596
rect 36596 22584 36602 22636
rect 36630 22584 36636 22636
rect 36688 22624 36694 22636
rect 37936 22633 37964 22664
rect 39482 22652 39488 22664
rect 39540 22652 39546 22704
rect 37277 22627 37335 22633
rect 37277 22624 37289 22627
rect 36688 22596 37289 22624
rect 36688 22584 36694 22596
rect 37277 22593 37289 22596
rect 37323 22593 37335 22627
rect 37277 22587 37335 22593
rect 37921 22627 37979 22633
rect 37921 22593 37933 22627
rect 37967 22593 37979 22627
rect 38654 22624 38660 22636
rect 38615 22596 38660 22624
rect 37921 22587 37979 22593
rect 38654 22584 38660 22596
rect 38712 22584 38718 22636
rect 39684 22633 39712 22732
rect 39853 22729 39865 22763
rect 39899 22760 39911 22763
rect 40034 22760 40040 22772
rect 39899 22732 40040 22760
rect 39899 22729 39911 22732
rect 39853 22723 39911 22729
rect 40034 22720 40040 22732
rect 40092 22720 40098 22772
rect 40770 22720 40776 22772
rect 40828 22760 40834 22772
rect 41049 22763 41107 22769
rect 41049 22760 41061 22763
rect 40828 22732 41061 22760
rect 40828 22720 40834 22732
rect 41049 22729 41061 22732
rect 41095 22729 41107 22763
rect 41049 22723 41107 22729
rect 41138 22720 41144 22772
rect 41196 22760 41202 22772
rect 41196 22732 47624 22760
rect 41196 22720 41202 22732
rect 39942 22652 39948 22704
rect 40000 22692 40006 22704
rect 40000 22664 40724 22692
rect 40000 22652 40006 22664
rect 39301 22627 39359 22633
rect 39301 22593 39313 22627
rect 39347 22593 39359 22627
rect 39301 22587 39359 22593
rect 39577 22627 39635 22633
rect 39577 22593 39589 22627
rect 39623 22593 39635 22627
rect 39577 22587 39635 22593
rect 39669 22627 39727 22633
rect 39669 22593 39681 22627
rect 39715 22624 39727 22627
rect 40126 22624 40132 22636
rect 39715 22596 40132 22624
rect 39715 22593 39727 22596
rect 39669 22587 39727 22593
rect 32306 22516 32312 22568
rect 32364 22556 32370 22568
rect 33045 22559 33103 22565
rect 33045 22556 33057 22559
rect 32364 22528 33057 22556
rect 32364 22516 32370 22528
rect 33045 22525 33057 22528
rect 33091 22525 33103 22559
rect 33045 22519 33103 22525
rect 37369 22491 37427 22497
rect 37369 22457 37381 22491
rect 37415 22488 37427 22491
rect 39316 22488 39344 22587
rect 39592 22556 39620 22587
rect 40126 22584 40132 22596
rect 40184 22584 40190 22636
rect 40310 22624 40316 22636
rect 40271 22596 40316 22624
rect 40310 22584 40316 22596
rect 40368 22584 40374 22636
rect 40402 22584 40408 22636
rect 40460 22624 40466 22636
rect 40696 22633 40724 22664
rect 45094 22652 45100 22704
rect 45152 22692 45158 22704
rect 45370 22692 45376 22704
rect 45152 22664 45376 22692
rect 45152 22652 45158 22664
rect 45370 22652 45376 22664
rect 45428 22692 45434 22704
rect 45465 22695 45523 22701
rect 45465 22692 45477 22695
rect 45428 22664 45477 22692
rect 45428 22652 45434 22664
rect 45465 22661 45477 22664
rect 45511 22661 45523 22695
rect 45465 22655 45523 22661
rect 40497 22627 40555 22633
rect 40497 22624 40509 22627
rect 40460 22596 40509 22624
rect 40460 22584 40466 22596
rect 40497 22593 40509 22596
rect 40543 22593 40555 22627
rect 40497 22587 40555 22593
rect 40681 22627 40739 22633
rect 40681 22593 40693 22627
rect 40727 22593 40739 22627
rect 40681 22587 40739 22593
rect 40865 22627 40923 22633
rect 40865 22593 40877 22627
rect 40911 22593 40923 22627
rect 40865 22587 40923 22593
rect 39758 22556 39764 22568
rect 39592 22528 39764 22556
rect 39758 22516 39764 22528
rect 39816 22516 39822 22568
rect 40586 22556 40592 22568
rect 40547 22528 40592 22556
rect 40586 22516 40592 22528
rect 40644 22516 40650 22568
rect 40880 22488 40908 22587
rect 42058 22584 42064 22636
rect 42116 22624 42122 22636
rect 42426 22624 42432 22636
rect 42116 22596 42432 22624
rect 42116 22584 42122 22596
rect 42426 22584 42432 22596
rect 42484 22584 42490 22636
rect 42518 22584 42524 22636
rect 42576 22624 42582 22636
rect 42685 22627 42743 22633
rect 42685 22624 42697 22627
rect 42576 22596 42697 22624
rect 42576 22584 42582 22596
rect 42685 22593 42697 22596
rect 42731 22593 42743 22627
rect 42685 22587 42743 22593
rect 45002 22584 45008 22636
rect 45060 22624 45066 22636
rect 47596 22633 47624 22732
rect 45281 22627 45339 22633
rect 45281 22624 45293 22627
rect 45060 22596 45293 22624
rect 45060 22584 45066 22596
rect 45281 22593 45293 22596
rect 45327 22593 45339 22627
rect 45281 22587 45339 22593
rect 47581 22627 47639 22633
rect 47581 22593 47593 22627
rect 47627 22593 47639 22627
rect 47581 22587 47639 22593
rect 41506 22488 41512 22500
rect 37415 22460 39252 22488
rect 39316 22460 41512 22488
rect 37415 22457 37427 22460
rect 37369 22451 37427 22457
rect 24302 22380 24308 22432
rect 24360 22420 24366 22432
rect 24397 22423 24455 22429
rect 24397 22420 24409 22423
rect 24360 22392 24409 22420
rect 24360 22380 24366 22392
rect 24397 22389 24409 22392
rect 24443 22389 24455 22423
rect 24397 22383 24455 22389
rect 31202 22380 31208 22432
rect 31260 22420 31266 22432
rect 31389 22423 31447 22429
rect 31389 22420 31401 22423
rect 31260 22392 31401 22420
rect 31260 22380 31266 22392
rect 31389 22389 31401 22392
rect 31435 22389 31447 22423
rect 31389 22383 31447 22389
rect 35897 22423 35955 22429
rect 35897 22389 35909 22423
rect 35943 22420 35955 22423
rect 36078 22420 36084 22432
rect 35943 22392 36084 22420
rect 35943 22389 35955 22392
rect 35897 22383 35955 22389
rect 36078 22380 36084 22392
rect 36136 22380 36142 22432
rect 38749 22423 38807 22429
rect 38749 22389 38761 22423
rect 38795 22420 38807 22423
rect 39114 22420 39120 22432
rect 38795 22392 39120 22420
rect 38795 22389 38807 22392
rect 38749 22383 38807 22389
rect 39114 22380 39120 22392
rect 39172 22380 39178 22432
rect 39224 22420 39252 22460
rect 41506 22448 41512 22460
rect 41564 22448 41570 22500
rect 40402 22420 40408 22432
rect 39224 22392 40408 22420
rect 40402 22380 40408 22392
rect 40460 22380 40466 22432
rect 43809 22423 43867 22429
rect 43809 22389 43821 22423
rect 43855 22420 43867 22423
rect 44174 22420 44180 22432
rect 43855 22392 44180 22420
rect 43855 22389 43867 22392
rect 43809 22383 43867 22389
rect 44174 22380 44180 22392
rect 44232 22380 44238 22432
rect 45646 22420 45652 22432
rect 45607 22392 45652 22420
rect 45646 22380 45652 22392
rect 45704 22380 45710 22432
rect 47026 22420 47032 22432
rect 46987 22392 47032 22420
rect 47026 22380 47032 22392
rect 47084 22380 47090 22432
rect 47670 22420 47676 22432
rect 47631 22392 47676 22420
rect 47670 22380 47676 22392
rect 47728 22380 47734 22432
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 25774 22216 25780 22228
rect 25735 22188 25780 22216
rect 25774 22176 25780 22188
rect 25832 22176 25838 22228
rect 26418 22216 26424 22228
rect 26379 22188 26424 22216
rect 26418 22176 26424 22188
rect 26476 22216 26482 22228
rect 26970 22216 26976 22228
rect 26476 22188 26976 22216
rect 26476 22176 26482 22188
rect 26970 22176 26976 22188
rect 27028 22176 27034 22228
rect 29822 22176 29828 22228
rect 29880 22216 29886 22228
rect 30009 22219 30067 22225
rect 30009 22216 30021 22219
rect 29880 22188 30021 22216
rect 29880 22176 29886 22188
rect 30009 22185 30021 22188
rect 30055 22185 30067 22219
rect 30374 22216 30380 22228
rect 30287 22188 30380 22216
rect 30009 22179 30067 22185
rect 30374 22176 30380 22188
rect 30432 22216 30438 22228
rect 31110 22216 31116 22228
rect 30432 22188 31116 22216
rect 30432 22176 30438 22188
rect 31110 22176 31116 22188
rect 31168 22176 31174 22228
rect 39114 22176 39120 22228
rect 39172 22216 39178 22228
rect 39850 22216 39856 22228
rect 39172 22188 39856 22216
rect 39172 22176 39178 22188
rect 39850 22176 39856 22188
rect 39908 22176 39914 22228
rect 40310 22176 40316 22228
rect 40368 22216 40374 22228
rect 40589 22219 40647 22225
rect 40589 22216 40601 22219
rect 40368 22188 40601 22216
rect 40368 22176 40374 22188
rect 40589 22185 40601 22188
rect 40635 22185 40647 22219
rect 40589 22179 40647 22185
rect 42429 22219 42487 22225
rect 42429 22185 42441 22219
rect 42475 22216 42487 22219
rect 42518 22216 42524 22228
rect 42475 22188 42524 22216
rect 42475 22185 42487 22188
rect 42429 22179 42487 22185
rect 42518 22176 42524 22188
rect 42576 22176 42582 22228
rect 17218 22108 17224 22160
rect 17276 22148 17282 22160
rect 17862 22148 17868 22160
rect 17276 22120 17868 22148
rect 17276 22108 17282 22120
rect 17862 22108 17868 22120
rect 17920 22108 17926 22160
rect 30466 22108 30472 22160
rect 30524 22108 30530 22160
rect 27341 22083 27399 22089
rect 27341 22049 27353 22083
rect 27387 22080 27399 22083
rect 27614 22080 27620 22092
rect 27387 22052 27620 22080
rect 27387 22049 27399 22052
rect 27341 22043 27399 22049
rect 27614 22040 27620 22052
rect 27672 22080 27678 22092
rect 28350 22080 28356 22092
rect 27672 22052 28356 22080
rect 27672 22040 27678 22052
rect 28350 22040 28356 22052
rect 28408 22080 28414 22092
rect 29362 22080 29368 22092
rect 28408 22052 29368 22080
rect 28408 22040 28414 22052
rect 29362 22040 29368 22052
rect 29420 22040 29426 22092
rect 30484 22080 30512 22108
rect 31018 22080 31024 22092
rect 30208 22052 30512 22080
rect 30979 22052 31024 22080
rect 2038 21972 2044 22024
rect 2096 22012 2102 22024
rect 2317 22015 2375 22021
rect 2317 22012 2329 22015
rect 2096 21984 2329 22012
rect 2096 21972 2102 21984
rect 2317 21981 2329 21984
rect 2363 21981 2375 22015
rect 2317 21975 2375 21981
rect 24397 22015 24455 22021
rect 24397 21981 24409 22015
rect 24443 22012 24455 22015
rect 27065 22015 27123 22021
rect 24443 21984 24900 22012
rect 24443 21981 24455 21984
rect 24397 21975 24455 21981
rect 24872 21956 24900 21984
rect 27065 21981 27077 22015
rect 27111 21981 27123 22015
rect 27065 21975 27123 21981
rect 24664 21947 24722 21953
rect 24664 21913 24676 21947
rect 24710 21944 24722 21947
rect 24762 21944 24768 21956
rect 24710 21916 24768 21944
rect 24710 21913 24722 21916
rect 24664 21907 24722 21913
rect 24762 21904 24768 21916
rect 24820 21904 24826 21956
rect 24854 21904 24860 21956
rect 24912 21904 24918 21956
rect 25774 21904 25780 21956
rect 25832 21944 25838 21956
rect 26237 21947 26295 21953
rect 26237 21944 26249 21947
rect 25832 21916 26249 21944
rect 25832 21904 25838 21916
rect 26237 21913 26249 21916
rect 26283 21944 26295 21947
rect 27080 21944 27108 21975
rect 27154 21972 27160 22024
rect 27212 22012 27218 22024
rect 30208 22021 30236 22052
rect 31018 22040 31024 22052
rect 31076 22040 31082 22092
rect 31110 22040 31116 22092
rect 31168 22080 31174 22092
rect 31297 22083 31355 22089
rect 31297 22080 31309 22083
rect 31168 22052 31309 22080
rect 31168 22040 31174 22052
rect 31297 22049 31309 22052
rect 31343 22049 31355 22083
rect 31297 22043 31355 22049
rect 31754 22040 31760 22092
rect 31812 22080 31818 22092
rect 32582 22080 32588 22092
rect 31812 22052 32588 22080
rect 31812 22040 31818 22052
rect 32582 22040 32588 22052
rect 32640 22040 32646 22092
rect 35434 22040 35440 22092
rect 35492 22080 35498 22092
rect 35805 22083 35863 22089
rect 35805 22080 35817 22083
rect 35492 22052 35817 22080
rect 35492 22040 35498 22052
rect 35805 22049 35817 22052
rect 35851 22049 35863 22083
rect 41414 22080 41420 22092
rect 35805 22043 35863 22049
rect 39776 22052 41420 22080
rect 30193 22015 30251 22021
rect 27212 21984 27257 22012
rect 27212 21972 27218 21984
rect 30193 21981 30205 22015
rect 30239 21981 30251 22015
rect 30193 21975 30251 21981
rect 30469 22015 30527 22021
rect 30469 21981 30481 22015
rect 30515 22012 30527 22015
rect 30558 22012 30564 22024
rect 30515 21984 30564 22012
rect 30515 21981 30527 21984
rect 30469 21975 30527 21981
rect 30558 21972 30564 21984
rect 30616 22012 30622 22024
rect 31202 22012 31208 22024
rect 30616 21984 31208 22012
rect 30616 21972 30622 21984
rect 31202 21972 31208 21984
rect 31260 21972 31266 22024
rect 32309 22015 32367 22021
rect 32309 21981 32321 22015
rect 32355 21981 32367 22015
rect 32309 21975 32367 21981
rect 38933 22015 38991 22021
rect 38933 21981 38945 22015
rect 38979 22012 38991 22015
rect 39574 22012 39580 22024
rect 38979 21984 39580 22012
rect 38979 21981 38991 21984
rect 38933 21975 38991 21981
rect 32324 21944 32352 21975
rect 39574 21972 39580 21984
rect 39632 21972 39638 22024
rect 34606 21944 34612 21956
rect 26283 21916 27108 21944
rect 27172 21916 34612 21944
rect 26283 21913 26295 21916
rect 26237 21907 26295 21913
rect 26418 21836 26424 21888
rect 26476 21885 26482 21888
rect 26476 21879 26495 21885
rect 26483 21845 26495 21879
rect 26602 21876 26608 21888
rect 26563 21848 26608 21876
rect 26476 21839 26495 21845
rect 26476 21836 26482 21839
rect 26602 21836 26608 21848
rect 26660 21836 26666 21888
rect 26694 21836 26700 21888
rect 26752 21876 26758 21888
rect 27172 21876 27200 21916
rect 34606 21904 34612 21916
rect 34664 21904 34670 21956
rect 35894 21904 35900 21956
rect 35952 21944 35958 21956
rect 36050 21947 36108 21953
rect 36050 21944 36062 21947
rect 35952 21916 36062 21944
rect 35952 21904 35958 21916
rect 36050 21913 36062 21916
rect 36096 21913 36108 21947
rect 36050 21907 36108 21913
rect 39117 21947 39175 21953
rect 39117 21913 39129 21947
rect 39163 21944 39175 21947
rect 39776 21944 39804 22052
rect 41414 22040 41420 22052
rect 41472 22080 41478 22092
rect 44174 22080 44180 22092
rect 41472 22052 44180 22080
rect 41472 22040 41478 22052
rect 39942 22012 39948 22024
rect 39903 21984 39948 22012
rect 39942 21972 39948 21984
rect 40000 21972 40006 22024
rect 40034 21972 40040 22024
rect 40092 22012 40098 22024
rect 40092 21984 40137 22012
rect 40092 21972 40098 21984
rect 40402 21972 40408 22024
rect 40460 22021 40466 22024
rect 40460 22012 40468 22021
rect 40460 21984 40505 22012
rect 40460 21975 40468 21984
rect 40460 21972 40466 21975
rect 40678 21972 40684 22024
rect 40736 22012 40742 22024
rect 41693 22015 41751 22021
rect 41693 22012 41705 22015
rect 40736 21984 41705 22012
rect 40736 21972 40742 21984
rect 41693 21981 41705 21984
rect 41739 21981 41751 22015
rect 41693 21975 41751 21981
rect 41782 21972 41788 22024
rect 41840 22012 41846 22024
rect 41877 22015 41935 22021
rect 41877 22012 41889 22015
rect 41840 21984 41889 22012
rect 41840 21972 41846 21984
rect 41877 21981 41889 21984
rect 41923 21981 41935 22015
rect 41969 22015 42027 22021
rect 41969 22002 41981 22015
rect 42015 22002 42027 22015
rect 42061 22015 42119 22021
rect 41877 21975 41935 21981
rect 39163 21916 39804 21944
rect 39163 21913 39175 21916
rect 39117 21907 39175 21913
rect 39850 21904 39856 21956
rect 39908 21944 39914 21956
rect 40221 21947 40279 21953
rect 40221 21944 40233 21947
rect 39908 21916 40233 21944
rect 39908 21904 39914 21916
rect 40221 21913 40233 21916
rect 40267 21913 40279 21947
rect 40221 21907 40279 21913
rect 40313 21947 40371 21953
rect 40313 21913 40325 21947
rect 40359 21944 40371 21947
rect 40586 21944 40592 21956
rect 40359 21916 40592 21944
rect 40359 21913 40371 21916
rect 40313 21907 40371 21913
rect 40586 21904 40592 21916
rect 40644 21904 40650 21956
rect 41966 21950 41972 22002
rect 42024 21950 42030 22002
rect 42061 21981 42073 22015
rect 42107 22012 42119 22015
rect 42150 22012 42156 22024
rect 42107 21984 42156 22012
rect 42107 21981 42119 21984
rect 42061 21975 42119 21981
rect 42150 21972 42156 21984
rect 42208 21972 42214 22024
rect 42260 22021 42288 22052
rect 44174 22040 44180 22052
rect 44232 22040 44238 22092
rect 45002 22040 45008 22092
rect 45060 22080 45066 22092
rect 45281 22083 45339 22089
rect 45281 22080 45293 22083
rect 45060 22052 45293 22080
rect 45060 22040 45066 22052
rect 45281 22049 45293 22052
rect 45327 22049 45339 22083
rect 45281 22043 45339 22049
rect 46293 22083 46351 22089
rect 46293 22049 46305 22083
rect 46339 22080 46351 22083
rect 47026 22080 47032 22092
rect 46339 22052 47032 22080
rect 46339 22049 46351 22052
rect 46293 22043 46351 22049
rect 47026 22040 47032 22052
rect 47084 22040 47090 22092
rect 48130 22080 48136 22092
rect 48091 22052 48136 22080
rect 48130 22040 48136 22052
rect 48188 22040 48194 22092
rect 42245 22015 42303 22021
rect 42245 21981 42257 22015
rect 42291 21981 42303 22015
rect 42245 21975 42303 21981
rect 42889 22015 42947 22021
rect 42889 21981 42901 22015
rect 42935 22012 42947 22015
rect 42978 22012 42984 22024
rect 42935 21984 42984 22012
rect 42935 21981 42947 21984
rect 42889 21975 42947 21981
rect 42978 21972 42984 21984
rect 43036 21972 43042 22024
rect 43073 22015 43131 22021
rect 43073 21981 43085 22015
rect 43119 21981 43131 22015
rect 43073 21975 43131 21981
rect 42702 21904 42708 21956
rect 42760 21944 42766 21956
rect 43088 21944 43116 21975
rect 44542 21972 44548 22024
rect 44600 22012 44606 22024
rect 45189 22015 45247 22021
rect 45189 22012 45201 22015
rect 44600 21984 45201 22012
rect 44600 21972 44606 21984
rect 45189 21981 45201 21984
rect 45235 21981 45247 22015
rect 45370 22012 45376 22024
rect 45331 21984 45376 22012
rect 45189 21975 45247 21981
rect 45370 21972 45376 21984
rect 45428 21972 45434 22024
rect 45462 21972 45468 22024
rect 45520 22012 45526 22024
rect 45520 21984 45565 22012
rect 45520 21972 45526 21984
rect 44726 21944 44732 21956
rect 42760 21916 44732 21944
rect 42760 21904 42766 21916
rect 44726 21904 44732 21916
rect 44784 21904 44790 21956
rect 46477 21947 46535 21953
rect 46477 21913 46489 21947
rect 46523 21944 46535 21947
rect 47670 21944 47676 21956
rect 46523 21916 47676 21944
rect 46523 21913 46535 21916
rect 46477 21907 46535 21913
rect 47670 21904 47676 21916
rect 47728 21904 47734 21956
rect 27338 21876 27344 21888
rect 26752 21848 27200 21876
rect 27299 21848 27344 21876
rect 26752 21836 26758 21848
rect 27338 21836 27344 21848
rect 27396 21836 27402 21888
rect 37182 21876 37188 21888
rect 37143 21848 37188 21876
rect 37182 21836 37188 21848
rect 37240 21836 37246 21888
rect 39301 21879 39359 21885
rect 39301 21845 39313 21879
rect 39347 21876 39359 21879
rect 39482 21876 39488 21888
rect 39347 21848 39488 21876
rect 39347 21845 39359 21848
rect 39301 21839 39359 21845
rect 39482 21836 39488 21848
rect 39540 21836 39546 21888
rect 40604 21876 40632 21904
rect 42610 21876 42616 21888
rect 40604 21848 42616 21876
rect 42610 21836 42616 21848
rect 42668 21836 42674 21888
rect 42978 21876 42984 21888
rect 42939 21848 42984 21876
rect 42978 21836 42984 21848
rect 43036 21836 43042 21888
rect 44266 21836 44272 21888
rect 44324 21876 44330 21888
rect 45005 21879 45063 21885
rect 45005 21876 45017 21879
rect 44324 21848 45017 21876
rect 44324 21836 44330 21848
rect 45005 21845 45017 21848
rect 45051 21845 45063 21879
rect 45005 21839 45063 21845
rect 45278 21836 45284 21888
rect 45336 21876 45342 21888
rect 45554 21876 45560 21888
rect 45336 21848 45560 21876
rect 45336 21836 45342 21848
rect 45554 21836 45560 21848
rect 45612 21836 45618 21888
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 25133 21675 25191 21681
rect 25133 21672 25145 21675
rect 24820 21644 25145 21672
rect 24820 21632 24826 21644
rect 25133 21641 25145 21644
rect 25179 21641 25191 21675
rect 25133 21635 25191 21641
rect 28810 21632 28816 21684
rect 28868 21632 28874 21684
rect 30374 21632 30380 21684
rect 30432 21681 30438 21684
rect 30432 21675 30451 21681
rect 30439 21641 30451 21675
rect 30432 21635 30451 21641
rect 30432 21632 30438 21635
rect 35894 21632 35900 21684
rect 35952 21672 35958 21684
rect 35952 21644 35997 21672
rect 35952 21632 35958 21644
rect 39942 21632 39948 21684
rect 40000 21672 40006 21684
rect 40221 21675 40279 21681
rect 40221 21672 40233 21675
rect 40000 21644 40233 21672
rect 40000 21632 40006 21644
rect 40221 21641 40233 21644
rect 40267 21641 40279 21675
rect 40221 21635 40279 21641
rect 41877 21675 41935 21681
rect 41877 21641 41889 21675
rect 41923 21672 41935 21675
rect 41966 21672 41972 21684
rect 41923 21644 41972 21672
rect 41923 21641 41935 21644
rect 41877 21635 41935 21641
rect 41966 21632 41972 21644
rect 42024 21632 42030 21684
rect 42978 21672 42984 21684
rect 42939 21644 42984 21672
rect 42978 21632 42984 21644
rect 43036 21632 43042 21684
rect 44910 21632 44916 21684
rect 44968 21672 44974 21684
rect 45005 21675 45063 21681
rect 45005 21672 45017 21675
rect 44968 21644 45017 21672
rect 44968 21632 44974 21644
rect 45005 21641 45017 21644
rect 45051 21672 45063 21675
rect 45278 21672 45284 21684
rect 45051 21644 45284 21672
rect 45051 21641 45063 21644
rect 45005 21635 45063 21641
rect 45278 21632 45284 21644
rect 45336 21632 45342 21684
rect 27338 21604 27344 21616
rect 25056 21576 27344 21604
rect 2038 21536 2044 21548
rect 1999 21508 2044 21536
rect 2038 21496 2044 21508
rect 2096 21496 2102 21548
rect 24302 21536 24308 21548
rect 24263 21508 24308 21536
rect 24302 21496 24308 21508
rect 24360 21496 24366 21548
rect 25056 21545 25084 21576
rect 27338 21564 27344 21576
rect 27396 21564 27402 21616
rect 28828 21604 28856 21632
rect 27908 21576 28856 21604
rect 30193 21607 30251 21613
rect 25041 21539 25099 21545
rect 25041 21505 25053 21539
rect 25087 21505 25099 21539
rect 25041 21499 25099 21505
rect 25225 21539 25283 21545
rect 25225 21505 25237 21539
rect 25271 21536 25283 21539
rect 26602 21536 26608 21548
rect 25271 21508 26608 21536
rect 25271 21505 25283 21508
rect 25225 21499 25283 21505
rect 2225 21471 2283 21477
rect 2225 21437 2237 21471
rect 2271 21468 2283 21471
rect 2406 21468 2412 21480
rect 2271 21440 2412 21468
rect 2271 21437 2283 21440
rect 2225 21431 2283 21437
rect 2406 21428 2412 21440
rect 2464 21428 2470 21480
rect 2774 21468 2780 21480
rect 2735 21440 2780 21468
rect 2774 21428 2780 21440
rect 2832 21428 2838 21480
rect 24578 21468 24584 21480
rect 24539 21440 24584 21468
rect 24578 21428 24584 21440
rect 24636 21428 24642 21480
rect 2866 21360 2872 21412
rect 2924 21400 2930 21412
rect 16758 21400 16764 21412
rect 2924 21372 16764 21400
rect 2924 21360 2930 21372
rect 16758 21360 16764 21372
rect 16816 21360 16822 21412
rect 24489 21403 24547 21409
rect 24489 21369 24501 21403
rect 24535 21400 24547 21403
rect 24670 21400 24676 21412
rect 24535 21372 24676 21400
rect 24535 21369 24547 21372
rect 24489 21363 24547 21369
rect 24670 21360 24676 21372
rect 24728 21400 24734 21412
rect 25240 21400 25268 21499
rect 26602 21496 26608 21508
rect 26660 21496 26666 21548
rect 27908 21545 27936 21576
rect 30193 21573 30205 21607
rect 30239 21604 30251 21607
rect 30558 21604 30564 21616
rect 30239 21576 30564 21604
rect 30239 21573 30251 21576
rect 30193 21567 30251 21573
rect 30558 21564 30564 21576
rect 30616 21564 30622 21616
rect 30650 21564 30656 21616
rect 30708 21604 30714 21616
rect 31021 21607 31079 21613
rect 31021 21604 31033 21607
rect 30708 21576 31033 21604
rect 30708 21564 30714 21576
rect 31021 21573 31033 21576
rect 31067 21573 31079 21607
rect 31021 21567 31079 21573
rect 31110 21564 31116 21616
rect 31168 21604 31174 21616
rect 42702 21604 42708 21616
rect 31168 21576 31340 21604
rect 31168 21564 31174 21576
rect 27157 21539 27215 21545
rect 27157 21536 27169 21539
rect 26896 21508 27169 21536
rect 26418 21428 26424 21480
rect 26476 21468 26482 21480
rect 26896 21468 26924 21508
rect 27157 21505 27169 21508
rect 27203 21505 27215 21539
rect 27157 21499 27215 21505
rect 27893 21539 27951 21545
rect 27893 21505 27905 21539
rect 27939 21505 27951 21539
rect 27893 21499 27951 21505
rect 27985 21539 28043 21545
rect 27985 21505 27997 21539
rect 28031 21536 28043 21539
rect 28258 21536 28264 21548
rect 28031 21508 28264 21536
rect 28031 21505 28043 21508
rect 27985 21499 28043 21505
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 28442 21496 28448 21548
rect 28500 21536 28506 21548
rect 28629 21539 28687 21545
rect 28629 21536 28641 21539
rect 28500 21508 28641 21536
rect 28500 21496 28506 21508
rect 28629 21505 28641 21508
rect 28675 21505 28687 21539
rect 28629 21499 28687 21505
rect 28813 21539 28871 21545
rect 28813 21505 28825 21539
rect 28859 21505 28871 21539
rect 31202 21536 31208 21548
rect 31163 21508 31208 21536
rect 28813 21499 28871 21505
rect 26476 21440 26924 21468
rect 26476 21428 26482 21440
rect 26970 21428 26976 21480
rect 27028 21468 27034 21480
rect 28828 21468 28856 21499
rect 31202 21496 31208 21508
rect 31260 21496 31266 21548
rect 31312 21545 31340 21576
rect 38856 21576 42708 21604
rect 38856 21548 38884 21576
rect 42702 21564 42708 21576
rect 42760 21564 42766 21616
rect 44542 21604 44548 21616
rect 42812 21576 44548 21604
rect 31297 21539 31355 21545
rect 31297 21505 31309 21539
rect 31343 21505 31355 21539
rect 34422 21536 34428 21548
rect 34383 21508 34428 21536
rect 31297 21499 31355 21505
rect 34422 21496 34428 21508
rect 34480 21496 34486 21548
rect 36078 21536 36084 21548
rect 36039 21508 36084 21536
rect 36078 21496 36084 21508
rect 36136 21496 36142 21548
rect 36265 21539 36323 21545
rect 36265 21505 36277 21539
rect 36311 21536 36323 21539
rect 36538 21536 36544 21548
rect 36311 21508 36544 21536
rect 36311 21505 36323 21508
rect 36265 21499 36323 21505
rect 36538 21496 36544 21508
rect 36596 21496 36602 21548
rect 38102 21496 38108 21548
rect 38160 21536 38166 21548
rect 38289 21539 38347 21545
rect 38289 21536 38301 21539
rect 38160 21508 38301 21536
rect 38160 21496 38166 21508
rect 38289 21505 38301 21508
rect 38335 21505 38347 21539
rect 38289 21499 38347 21505
rect 38473 21539 38531 21545
rect 38473 21505 38485 21539
rect 38519 21505 38531 21539
rect 38654 21536 38660 21548
rect 38615 21508 38660 21536
rect 38473 21499 38531 21505
rect 27028 21440 27073 21468
rect 28184 21440 28856 21468
rect 36357 21471 36415 21477
rect 27028 21428 27034 21440
rect 24728 21372 25268 21400
rect 24728 21360 24734 21372
rect 24118 21332 24124 21344
rect 24079 21304 24124 21332
rect 24118 21292 24124 21304
rect 24176 21292 24182 21344
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 27154 21332 27160 21344
rect 26292 21304 27160 21332
rect 26292 21292 26298 21304
rect 27154 21292 27160 21304
rect 27212 21332 27218 21344
rect 27341 21335 27399 21341
rect 27341 21332 27353 21335
rect 27212 21304 27353 21332
rect 27212 21292 27218 21304
rect 27341 21301 27353 21304
rect 27387 21301 27399 21335
rect 27341 21295 27399 21301
rect 27982 21292 27988 21344
rect 28040 21332 28046 21344
rect 28184 21341 28212 21440
rect 36357 21437 36369 21471
rect 36403 21468 36415 21471
rect 37182 21468 37188 21480
rect 36403 21440 37188 21468
rect 36403 21437 36415 21440
rect 36357 21431 36415 21437
rect 37182 21428 37188 21440
rect 37240 21428 37246 21480
rect 30282 21360 30288 21412
rect 30340 21400 30346 21412
rect 30561 21403 30619 21409
rect 30561 21400 30573 21403
rect 30340 21372 30573 21400
rect 30340 21360 30346 21372
rect 30561 21369 30573 21372
rect 30607 21369 30619 21403
rect 30561 21363 30619 21369
rect 33870 21360 33876 21412
rect 33928 21400 33934 21412
rect 34517 21403 34575 21409
rect 34517 21400 34529 21403
rect 33928 21372 34529 21400
rect 33928 21360 33934 21372
rect 34517 21369 34529 21372
rect 34563 21400 34575 21403
rect 37918 21400 37924 21412
rect 34563 21372 37924 21400
rect 34563 21369 34575 21372
rect 34517 21363 34575 21369
rect 37918 21360 37924 21372
rect 37976 21400 37982 21412
rect 38488 21400 38516 21499
rect 38654 21496 38660 21508
rect 38712 21496 38718 21548
rect 38838 21536 38844 21548
rect 38799 21508 38844 21536
rect 38838 21496 38844 21508
rect 38896 21496 38902 21548
rect 39482 21536 39488 21548
rect 39443 21508 39488 21536
rect 39482 21496 39488 21508
rect 39540 21496 39546 21548
rect 39669 21539 39727 21545
rect 39669 21505 39681 21539
rect 39715 21505 39727 21539
rect 39850 21536 39856 21548
rect 39811 21508 39856 21536
rect 39669 21499 39727 21505
rect 38562 21428 38568 21480
rect 38620 21468 38626 21480
rect 39025 21471 39083 21477
rect 38620 21440 38665 21468
rect 38620 21428 38626 21440
rect 39025 21437 39037 21471
rect 39071 21468 39083 21471
rect 39684 21468 39712 21499
rect 39850 21496 39856 21508
rect 39908 21496 39914 21548
rect 40034 21536 40040 21548
rect 39995 21508 40040 21536
rect 40034 21496 40040 21508
rect 40092 21496 40098 21548
rect 41693 21539 41751 21545
rect 41693 21505 41705 21539
rect 41739 21505 41751 21539
rect 41874 21536 41880 21548
rect 41835 21508 41880 21536
rect 41693 21499 41751 21505
rect 39071 21440 39712 21468
rect 39071 21437 39083 21440
rect 39025 21431 39083 21437
rect 39758 21428 39764 21480
rect 39816 21468 39822 21480
rect 41708 21468 41736 21499
rect 41874 21496 41880 21508
rect 41932 21496 41938 21548
rect 42812 21545 42840 21576
rect 44542 21564 44548 21576
rect 44600 21564 44606 21616
rect 44726 21564 44732 21616
rect 44784 21604 44790 21616
rect 44784 21576 46152 21604
rect 44784 21564 44790 21576
rect 42797 21539 42855 21545
rect 42797 21505 42809 21539
rect 42843 21536 42855 21539
rect 42886 21536 42892 21548
rect 42843 21508 42892 21536
rect 42843 21505 42855 21508
rect 42797 21499 42855 21505
rect 42886 21496 42892 21508
rect 42944 21496 42950 21548
rect 43070 21536 43076 21548
rect 43031 21508 43076 21536
rect 43070 21496 43076 21508
rect 43128 21496 43134 21548
rect 44174 21536 44180 21548
rect 44087 21508 44180 21536
rect 44174 21496 44180 21508
rect 44232 21536 44238 21548
rect 44910 21536 44916 21548
rect 44232 21508 44916 21536
rect 44232 21496 44238 21508
rect 44910 21496 44916 21508
rect 44968 21496 44974 21548
rect 45373 21539 45431 21545
rect 45373 21505 45385 21539
rect 45419 21536 45431 21539
rect 45646 21536 45652 21548
rect 45419 21508 45652 21536
rect 45419 21505 45431 21508
rect 45373 21499 45431 21505
rect 45646 21496 45652 21508
rect 45704 21496 45710 21548
rect 42613 21471 42671 21477
rect 42613 21468 42625 21471
rect 39816 21440 39861 21468
rect 41708 21440 42625 21468
rect 39816 21428 39822 21440
rect 42613 21437 42625 21440
rect 42659 21437 42671 21471
rect 42613 21431 42671 21437
rect 44269 21471 44327 21477
rect 44269 21437 44281 21471
rect 44315 21468 44327 21471
rect 44358 21468 44364 21480
rect 44315 21440 44364 21468
rect 44315 21437 44327 21440
rect 44269 21431 44327 21437
rect 44358 21428 44364 21440
rect 44416 21428 44422 21480
rect 44542 21468 44548 21480
rect 44503 21440 44548 21468
rect 44542 21428 44548 21440
rect 44600 21428 44606 21480
rect 45094 21428 45100 21480
rect 45152 21468 45158 21480
rect 45465 21471 45523 21477
rect 45465 21468 45477 21471
rect 45152 21440 45477 21468
rect 45152 21428 45158 21440
rect 45465 21437 45477 21440
rect 45511 21437 45523 21471
rect 46124 21468 46152 21576
rect 46201 21539 46259 21545
rect 46201 21505 46213 21539
rect 46247 21536 46259 21539
rect 47765 21539 47823 21545
rect 47765 21536 47777 21539
rect 46247 21508 47777 21536
rect 46247 21505 46259 21508
rect 46201 21499 46259 21505
rect 47765 21505 47777 21508
rect 47811 21536 47823 21539
rect 48130 21536 48136 21548
rect 47811 21508 48136 21536
rect 47811 21505 47823 21508
rect 47765 21499 47823 21505
rect 48130 21496 48136 21508
rect 48188 21496 48194 21548
rect 46477 21471 46535 21477
rect 46477 21468 46489 21471
rect 46124 21440 46489 21468
rect 45465 21431 45523 21437
rect 46477 21437 46489 21440
rect 46523 21437 46535 21471
rect 47670 21468 47676 21480
rect 47631 21440 47676 21468
rect 46477 21431 46535 21437
rect 47670 21428 47676 21440
rect 47728 21428 47734 21480
rect 48133 21403 48191 21409
rect 48133 21400 48145 21403
rect 37976 21372 38516 21400
rect 45020 21372 48145 21400
rect 37976 21360 37982 21372
rect 45020 21344 45048 21372
rect 48133 21369 48145 21372
rect 48179 21369 48191 21403
rect 48133 21363 48191 21369
rect 28169 21335 28227 21341
rect 28169 21332 28181 21335
rect 28040 21304 28181 21332
rect 28040 21292 28046 21304
rect 28169 21301 28181 21304
rect 28215 21301 28227 21335
rect 28626 21332 28632 21344
rect 28587 21304 28632 21332
rect 28169 21295 28227 21301
rect 28626 21292 28632 21304
rect 28684 21292 28690 21344
rect 30377 21335 30435 21341
rect 30377 21301 30389 21335
rect 30423 21332 30435 21335
rect 30650 21332 30656 21344
rect 30423 21304 30656 21332
rect 30423 21301 30435 21304
rect 30377 21295 30435 21301
rect 30650 21292 30656 21304
rect 30708 21292 30714 21344
rect 31018 21332 31024 21344
rect 30979 21304 31024 21332
rect 31018 21292 31024 21304
rect 31076 21292 31082 21344
rect 38562 21292 38568 21344
rect 38620 21332 38626 21344
rect 43254 21332 43260 21344
rect 38620 21304 43260 21332
rect 38620 21292 38626 21304
rect 43254 21292 43260 21304
rect 43312 21292 43318 21344
rect 45002 21292 45008 21344
rect 45060 21292 45066 21344
rect 45649 21335 45707 21341
rect 45649 21301 45661 21335
rect 45695 21332 45707 21335
rect 46106 21332 46112 21344
rect 45695 21304 46112 21332
rect 45695 21301 45707 21304
rect 45649 21295 45707 21301
rect 46106 21292 46112 21304
rect 46164 21292 46170 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 2406 21128 2412 21140
rect 2367 21100 2412 21128
rect 2406 21088 2412 21100
rect 2464 21088 2470 21140
rect 24578 21088 24584 21140
rect 24636 21128 24642 21140
rect 25777 21131 25835 21137
rect 25777 21128 25789 21131
rect 24636 21100 25789 21128
rect 24636 21088 24642 21100
rect 25777 21097 25789 21100
rect 25823 21097 25835 21131
rect 25777 21091 25835 21097
rect 26973 21131 27031 21137
rect 26973 21097 26985 21131
rect 27019 21128 27031 21131
rect 27982 21128 27988 21140
rect 27019 21100 27988 21128
rect 27019 21097 27031 21100
rect 26973 21091 27031 21097
rect 27982 21088 27988 21100
rect 28040 21088 28046 21140
rect 28810 21088 28816 21140
rect 28868 21128 28874 21140
rect 28997 21131 29055 21137
rect 28997 21128 29009 21131
rect 28868 21100 29009 21128
rect 28868 21088 28874 21100
rect 28997 21097 29009 21100
rect 29043 21097 29055 21131
rect 28997 21091 29055 21097
rect 31297 21131 31355 21137
rect 31297 21097 31309 21131
rect 31343 21128 31355 21131
rect 31570 21128 31576 21140
rect 31343 21100 31576 21128
rect 31343 21097 31355 21100
rect 31297 21091 31355 21097
rect 31570 21088 31576 21100
rect 31628 21088 31634 21140
rect 38102 21128 38108 21140
rect 38063 21100 38108 21128
rect 38102 21088 38108 21100
rect 38160 21088 38166 21140
rect 39758 21088 39764 21140
rect 39816 21128 39822 21140
rect 40405 21131 40463 21137
rect 40405 21128 40417 21131
rect 39816 21100 40417 21128
rect 39816 21088 39822 21100
rect 40405 21097 40417 21100
rect 40451 21097 40463 21131
rect 40405 21091 40463 21097
rect 42981 21131 43039 21137
rect 42981 21097 42993 21131
rect 43027 21128 43039 21131
rect 43070 21128 43076 21140
rect 43027 21100 43076 21128
rect 43027 21097 43039 21100
rect 42981 21091 43039 21097
rect 43070 21088 43076 21100
rect 43128 21128 43134 21140
rect 45094 21128 45100 21140
rect 43128 21100 45100 21128
rect 43128 21088 43134 21100
rect 45094 21088 45100 21100
rect 45152 21088 45158 21140
rect 45186 21088 45192 21140
rect 45244 21128 45250 21140
rect 47670 21128 47676 21140
rect 45244 21100 47676 21128
rect 45244 21088 45250 21100
rect 47670 21088 47676 21100
rect 47728 21088 47734 21140
rect 48130 21128 48136 21140
rect 48091 21100 48136 21128
rect 48130 21088 48136 21100
rect 48188 21088 48194 21140
rect 27614 21020 27620 21072
rect 27672 21020 27678 21072
rect 33318 21020 33324 21072
rect 33376 21060 33382 21072
rect 33689 21063 33747 21069
rect 33689 21060 33701 21063
rect 33376 21032 33701 21060
rect 33376 21020 33382 21032
rect 33689 21029 33701 21032
rect 33735 21029 33747 21063
rect 33689 21023 33747 21029
rect 39025 21063 39083 21069
rect 39025 21029 39037 21063
rect 39071 21060 39083 21063
rect 39114 21060 39120 21072
rect 39071 21032 39120 21060
rect 39071 21029 39083 21032
rect 39025 21023 39083 21029
rect 39114 21020 39120 21032
rect 39172 21020 39178 21072
rect 41782 21020 41788 21072
rect 41840 21060 41846 21072
rect 43165 21063 43223 21069
rect 43165 21060 43177 21063
rect 41840 21032 43177 21060
rect 41840 21020 41846 21032
rect 43165 21029 43177 21032
rect 43211 21029 43223 21063
rect 43165 21023 43223 21029
rect 44358 21020 44364 21072
rect 44416 21060 44422 21072
rect 44818 21060 44824 21072
rect 44416 21032 44824 21060
rect 44416 21020 44422 21032
rect 44818 21020 44824 21032
rect 44876 21060 44882 21072
rect 45204 21060 45232 21088
rect 44876 21032 45232 21060
rect 44876 21020 44882 21032
rect 27157 20995 27215 21001
rect 27157 20961 27169 20995
rect 27203 20992 27215 20995
rect 27632 20992 27660 21020
rect 27203 20964 27660 20992
rect 27203 20961 27215 20964
rect 27157 20955 27215 20961
rect 29546 20952 29552 21004
rect 29604 20992 29610 21004
rect 29914 20992 29920 21004
rect 29604 20964 29920 20992
rect 29604 20952 29610 20964
rect 29914 20952 29920 20964
rect 29972 20952 29978 21004
rect 31202 20952 31208 21004
rect 31260 20992 31266 21004
rect 31260 20964 31984 20992
rect 31260 20952 31266 20964
rect 2317 20927 2375 20933
rect 2317 20893 2329 20927
rect 2363 20924 2375 20927
rect 2866 20924 2872 20936
rect 2363 20896 2872 20924
rect 2363 20893 2375 20896
rect 2317 20887 2375 20893
rect 2866 20884 2872 20896
rect 2924 20884 2930 20936
rect 3142 20924 3148 20936
rect 3103 20896 3148 20924
rect 3142 20884 3148 20896
rect 3200 20884 3206 20936
rect 24397 20927 24455 20933
rect 24397 20893 24409 20927
rect 24443 20924 24455 20927
rect 24443 20896 24900 20924
rect 24443 20893 24455 20896
rect 24397 20887 24455 20893
rect 24872 20868 24900 20896
rect 26234 20884 26240 20936
rect 26292 20924 26298 20936
rect 26421 20927 26479 20933
rect 26292 20896 26337 20924
rect 26292 20884 26298 20896
rect 26421 20893 26433 20927
rect 26467 20924 26479 20927
rect 26694 20924 26700 20936
rect 26467 20896 26700 20924
rect 26467 20893 26479 20896
rect 26421 20887 26479 20893
rect 26694 20884 26700 20896
rect 26752 20884 26758 20936
rect 26881 20927 26939 20933
rect 26881 20893 26893 20927
rect 26927 20924 26939 20927
rect 27338 20924 27344 20936
rect 26927 20896 27344 20924
rect 26927 20893 26939 20896
rect 26881 20887 26939 20893
rect 27338 20884 27344 20896
rect 27396 20884 27402 20936
rect 27617 20927 27675 20933
rect 27617 20893 27629 20927
rect 27663 20924 27675 20927
rect 29564 20924 29592 20952
rect 31754 20924 31760 20936
rect 27663 20896 29592 20924
rect 31715 20896 31760 20924
rect 27663 20893 27675 20896
rect 27617 20887 27675 20893
rect 24118 20816 24124 20868
rect 24176 20856 24182 20868
rect 24642 20859 24700 20865
rect 24642 20856 24654 20859
rect 24176 20828 24654 20856
rect 24176 20816 24182 20828
rect 24642 20825 24654 20828
rect 24688 20825 24700 20859
rect 24642 20819 24700 20825
rect 24854 20816 24860 20868
rect 24912 20856 24918 20868
rect 27632 20856 27660 20887
rect 31754 20884 31760 20896
rect 31812 20884 31818 20936
rect 31956 20933 31984 20964
rect 34606 20952 34612 21004
rect 34664 20992 34670 21004
rect 38194 20992 38200 21004
rect 34664 20964 34928 20992
rect 34664 20952 34670 20964
rect 31941 20927 31999 20933
rect 31941 20893 31953 20927
rect 31987 20893 31999 20927
rect 33870 20924 33876 20936
rect 33831 20896 33876 20924
rect 31941 20887 31999 20893
rect 33870 20884 33876 20896
rect 33928 20884 33934 20936
rect 33965 20927 34023 20933
rect 33965 20893 33977 20927
rect 34011 20924 34023 20927
rect 34790 20924 34796 20936
rect 34011 20896 34796 20924
rect 34011 20893 34023 20896
rect 33965 20887 34023 20893
rect 34790 20884 34796 20896
rect 34848 20884 34854 20936
rect 34900 20933 34928 20964
rect 37844 20964 38200 20992
rect 34885 20927 34943 20933
rect 34885 20893 34897 20927
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 34974 20884 34980 20936
rect 35032 20924 35038 20936
rect 35161 20927 35219 20933
rect 35161 20924 35173 20927
rect 35032 20896 35173 20924
rect 35032 20884 35038 20896
rect 35161 20893 35173 20896
rect 35207 20893 35219 20927
rect 35618 20924 35624 20936
rect 35579 20896 35624 20924
rect 35161 20887 35219 20893
rect 35618 20884 35624 20896
rect 35676 20884 35682 20936
rect 37458 20924 37464 20936
rect 37419 20896 37464 20924
rect 37458 20884 37464 20896
rect 37516 20884 37522 20936
rect 37609 20927 37667 20933
rect 37609 20893 37621 20927
rect 37655 20924 37667 20927
rect 37844 20924 37872 20964
rect 38194 20952 38200 20964
rect 38252 20952 38258 21004
rect 38838 20952 38844 21004
rect 38896 20992 38902 21004
rect 38896 20964 39528 20992
rect 38896 20952 38902 20964
rect 37655 20896 37872 20924
rect 37655 20893 37667 20896
rect 37609 20887 37667 20893
rect 37918 20884 37924 20936
rect 37976 20933 37982 20936
rect 37976 20924 37984 20933
rect 39022 20924 39028 20936
rect 37976 20896 38021 20924
rect 38983 20896 39028 20924
rect 37976 20887 37984 20896
rect 37976 20884 37982 20887
rect 39022 20884 39028 20896
rect 39080 20884 39086 20936
rect 39298 20924 39304 20936
rect 39259 20896 39304 20924
rect 39298 20884 39304 20896
rect 39356 20884 39362 20936
rect 39500 20924 39528 20964
rect 39574 20952 39580 21004
rect 39632 20992 39638 21004
rect 39632 20964 40264 20992
rect 39632 20952 39638 20964
rect 40236 20933 40264 20964
rect 44726 20952 44732 21004
rect 44784 20992 44790 21004
rect 46750 20992 46756 21004
rect 44784 20964 45508 20992
rect 46711 20964 46756 20992
rect 44784 20952 44790 20964
rect 39853 20927 39911 20933
rect 39853 20924 39865 20927
rect 39500 20896 39865 20924
rect 39853 20893 39865 20896
rect 39899 20893 39911 20927
rect 39853 20887 39911 20893
rect 40221 20927 40279 20933
rect 40221 20893 40233 20927
rect 40267 20893 40279 20927
rect 40221 20887 40279 20893
rect 42978 20884 42984 20936
rect 43036 20884 43042 20936
rect 45002 20924 45008 20936
rect 44963 20896 45008 20924
rect 45002 20884 45008 20896
rect 45060 20884 45066 20936
rect 45189 20927 45247 20933
rect 45189 20893 45201 20927
rect 45235 20924 45247 20927
rect 45370 20924 45376 20936
rect 45235 20896 45376 20924
rect 45235 20893 45247 20896
rect 45189 20887 45247 20893
rect 45370 20884 45376 20896
rect 45428 20884 45434 20936
rect 45480 20924 45508 20964
rect 46750 20952 46756 20964
rect 46808 20952 46814 21004
rect 45879 20927 45937 20933
rect 45879 20924 45891 20927
rect 45480 20896 45891 20924
rect 45879 20893 45891 20896
rect 45925 20893 45937 20927
rect 46014 20924 46020 20936
rect 45975 20896 46020 20924
rect 45879 20887 45937 20893
rect 46014 20884 46020 20896
rect 46072 20884 46078 20936
rect 46106 20884 46112 20936
rect 46164 20924 46170 20936
rect 46164 20896 46209 20924
rect 46164 20884 46170 20896
rect 46290 20884 46296 20936
rect 46348 20924 46354 20936
rect 46348 20896 46393 20924
rect 46348 20884 46354 20896
rect 24912 20828 27660 20856
rect 27884 20859 27942 20865
rect 24912 20816 24918 20828
rect 27884 20825 27896 20859
rect 27930 20856 27942 20859
rect 28626 20856 28632 20868
rect 27930 20828 28632 20856
rect 27930 20825 27942 20828
rect 27884 20819 27942 20825
rect 28626 20816 28632 20828
rect 28684 20816 28690 20868
rect 30184 20859 30242 20865
rect 30184 20825 30196 20859
rect 30230 20856 30242 20859
rect 31849 20859 31907 20865
rect 31849 20856 31861 20859
rect 30230 20828 31861 20856
rect 30230 20825 30242 20828
rect 30184 20819 30242 20825
rect 31849 20825 31861 20828
rect 31895 20825 31907 20859
rect 31849 20819 31907 20825
rect 33689 20859 33747 20865
rect 33689 20825 33701 20859
rect 33735 20856 33747 20859
rect 34701 20859 34759 20865
rect 34701 20856 34713 20859
rect 33735 20828 34713 20856
rect 33735 20825 33747 20828
rect 33689 20819 33747 20825
rect 34701 20825 34713 20828
rect 34747 20825 34759 20859
rect 37734 20856 37740 20868
rect 37695 20828 37740 20856
rect 34701 20819 34759 20825
rect 37734 20816 37740 20828
rect 37792 20816 37798 20868
rect 37829 20859 37887 20865
rect 37829 20825 37841 20859
rect 37875 20856 37887 20859
rect 38562 20856 38568 20868
rect 37875 20828 38568 20856
rect 37875 20825 37887 20828
rect 37829 20819 37887 20825
rect 38562 20816 38568 20828
rect 38620 20816 38626 20868
rect 40037 20859 40095 20865
rect 40037 20856 40049 20859
rect 39132 20828 40049 20856
rect 26234 20748 26240 20800
rect 26292 20788 26298 20800
rect 26329 20791 26387 20797
rect 26329 20788 26341 20791
rect 26292 20760 26341 20788
rect 26292 20748 26298 20760
rect 26329 20757 26341 20760
rect 26375 20757 26387 20791
rect 26329 20751 26387 20757
rect 27062 20748 27068 20800
rect 27120 20788 27126 20800
rect 27157 20791 27215 20797
rect 27157 20788 27169 20791
rect 27120 20760 27169 20788
rect 27120 20748 27126 20760
rect 27157 20757 27169 20760
rect 27203 20757 27215 20791
rect 27157 20751 27215 20757
rect 34422 20748 34428 20800
rect 34480 20788 34486 20800
rect 35069 20791 35127 20797
rect 35069 20788 35081 20791
rect 34480 20760 35081 20788
rect 34480 20748 34486 20760
rect 35069 20757 35081 20760
rect 35115 20757 35127 20791
rect 35069 20751 35127 20757
rect 35713 20791 35771 20797
rect 35713 20757 35725 20791
rect 35759 20788 35771 20791
rect 38654 20788 38660 20800
rect 35759 20760 38660 20788
rect 35759 20757 35771 20760
rect 35713 20751 35771 20757
rect 38654 20748 38660 20760
rect 38712 20788 38718 20800
rect 39132 20788 39160 20828
rect 40037 20825 40049 20828
rect 40083 20825 40095 20859
rect 40037 20819 40095 20825
rect 40129 20859 40187 20865
rect 40129 20825 40141 20859
rect 40175 20856 40187 20859
rect 41414 20856 41420 20868
rect 40175 20828 41420 20856
rect 40175 20825 40187 20828
rect 40129 20819 40187 20825
rect 41414 20816 41420 20828
rect 41472 20816 41478 20868
rect 42797 20859 42855 20865
rect 42797 20825 42809 20859
rect 42843 20856 42855 20859
rect 42996 20856 43024 20884
rect 42843 20828 43024 20856
rect 45649 20859 45707 20865
rect 42843 20825 42855 20828
rect 42797 20819 42855 20825
rect 45649 20825 45661 20859
rect 45695 20856 45707 20859
rect 46998 20859 47056 20865
rect 46998 20856 47010 20859
rect 45695 20828 47010 20856
rect 45695 20825 45707 20828
rect 45649 20819 45707 20825
rect 46998 20825 47010 20828
rect 47044 20825 47056 20859
rect 46998 20819 47056 20825
rect 38712 20760 39160 20788
rect 39209 20791 39267 20797
rect 38712 20748 38718 20760
rect 39209 20757 39221 20791
rect 39255 20788 39267 20791
rect 39482 20788 39488 20800
rect 39255 20760 39488 20788
rect 39255 20757 39267 20760
rect 39209 20751 39267 20757
rect 39482 20748 39488 20760
rect 39540 20788 39546 20800
rect 42702 20788 42708 20800
rect 39540 20760 42708 20788
rect 39540 20748 39546 20760
rect 42702 20748 42708 20760
rect 42760 20748 42766 20800
rect 42886 20748 42892 20800
rect 42944 20788 42950 20800
rect 42997 20791 43055 20797
rect 42997 20788 43009 20791
rect 42944 20760 43009 20788
rect 42944 20748 42950 20760
rect 42997 20757 43009 20760
rect 43043 20757 43055 20791
rect 42997 20751 43055 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 28442 20584 28448 20596
rect 28403 20556 28448 20584
rect 28442 20544 28448 20556
rect 28500 20544 28506 20596
rect 30650 20544 30656 20596
rect 30708 20584 30714 20596
rect 31297 20587 31355 20593
rect 31297 20584 31309 20587
rect 30708 20556 31309 20584
rect 30708 20544 30714 20556
rect 31297 20553 31309 20556
rect 31343 20553 31355 20587
rect 34698 20584 34704 20596
rect 31297 20547 31355 20553
rect 33060 20556 34704 20584
rect 3142 20516 3148 20528
rect 2148 20488 3148 20516
rect 2148 20457 2176 20488
rect 3142 20476 3148 20488
rect 3200 20476 3206 20528
rect 27338 20516 27344 20528
rect 27299 20488 27344 20516
rect 27338 20476 27344 20488
rect 27396 20476 27402 20528
rect 27557 20519 27615 20525
rect 27557 20485 27569 20519
rect 27603 20516 27615 20519
rect 28258 20516 28264 20528
rect 27603 20488 28264 20516
rect 27603 20485 27615 20488
rect 27557 20479 27615 20485
rect 28258 20476 28264 20488
rect 28316 20476 28322 20528
rect 33060 20525 33088 20556
rect 34698 20544 34704 20556
rect 34756 20544 34762 20596
rect 34790 20544 34796 20596
rect 34848 20584 34854 20596
rect 35713 20587 35771 20593
rect 35713 20584 35725 20587
rect 34848 20556 35725 20584
rect 34848 20544 34854 20556
rect 35713 20553 35725 20556
rect 35759 20584 35771 20587
rect 37277 20587 37335 20593
rect 35759 20556 35894 20584
rect 35759 20553 35771 20556
rect 35713 20547 35771 20553
rect 33045 20519 33103 20525
rect 33045 20485 33057 20519
rect 33091 20485 33103 20519
rect 35434 20516 35440 20528
rect 33045 20479 33103 20485
rect 33796 20488 35440 20516
rect 2133 20451 2191 20457
rect 2133 20417 2145 20451
rect 2179 20417 2191 20451
rect 2133 20411 2191 20417
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 26234 20448 26240 20460
rect 26099 20420 26240 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 26234 20408 26240 20420
rect 26292 20408 26298 20460
rect 26326 20408 26332 20460
rect 26384 20448 26390 20460
rect 26970 20448 26976 20460
rect 26384 20420 26976 20448
rect 26384 20408 26390 20420
rect 26970 20408 26976 20420
rect 27028 20408 27034 20460
rect 28169 20451 28227 20457
rect 28169 20417 28181 20451
rect 28215 20448 28227 20451
rect 28810 20448 28816 20460
rect 28215 20420 28816 20448
rect 28215 20417 28227 20420
rect 28169 20411 28227 20417
rect 2317 20383 2375 20389
rect 2317 20349 2329 20383
rect 2363 20380 2375 20383
rect 2590 20380 2596 20392
rect 2363 20352 2596 20380
rect 2363 20349 2375 20352
rect 2317 20343 2375 20349
rect 2590 20340 2596 20352
rect 2648 20340 2654 20392
rect 2774 20380 2780 20392
rect 2735 20352 2780 20380
rect 2774 20340 2780 20352
rect 2832 20340 2838 20392
rect 26237 20315 26295 20321
rect 26237 20281 26249 20315
rect 26283 20312 26295 20315
rect 26418 20312 26424 20324
rect 26283 20284 26424 20312
rect 26283 20281 26295 20284
rect 26237 20275 26295 20281
rect 26418 20272 26424 20284
rect 26476 20312 26482 20324
rect 27246 20312 27252 20324
rect 26476 20284 27252 20312
rect 26476 20272 26482 20284
rect 27246 20272 27252 20284
rect 27304 20312 27310 20324
rect 27709 20315 27767 20321
rect 27709 20312 27721 20315
rect 27304 20284 27721 20312
rect 27304 20272 27310 20284
rect 27709 20281 27721 20284
rect 27755 20281 27767 20315
rect 28184 20312 28212 20411
rect 28810 20408 28816 20420
rect 28868 20408 28874 20460
rect 29914 20448 29920 20460
rect 29875 20420 29920 20448
rect 29914 20408 29920 20420
rect 29972 20408 29978 20460
rect 30190 20457 30196 20460
rect 30184 20411 30196 20457
rect 30248 20448 30254 20460
rect 33226 20448 33232 20460
rect 30248 20420 30284 20448
rect 33187 20420 33232 20448
rect 30190 20408 30196 20411
rect 30248 20408 30254 20420
rect 33226 20408 33232 20420
rect 33284 20408 33290 20460
rect 33321 20451 33379 20457
rect 33321 20417 33333 20451
rect 33367 20448 33379 20451
rect 33410 20448 33416 20460
rect 33367 20420 33416 20448
rect 33367 20417 33379 20420
rect 33321 20411 33379 20417
rect 33410 20408 33416 20420
rect 33468 20408 33474 20460
rect 33796 20457 33824 20488
rect 35434 20476 35440 20488
rect 35492 20476 35498 20528
rect 35866 20516 35894 20556
rect 37277 20553 37289 20587
rect 37323 20584 37335 20587
rect 37458 20584 37464 20596
rect 37323 20556 37464 20584
rect 37323 20553 37335 20556
rect 37277 20547 37335 20553
rect 37458 20544 37464 20556
rect 37516 20544 37522 20596
rect 37734 20584 37740 20596
rect 37660 20556 37740 20584
rect 37660 20516 37688 20556
rect 37734 20544 37740 20556
rect 37792 20544 37798 20596
rect 39298 20544 39304 20596
rect 39356 20584 39362 20596
rect 41690 20584 41696 20596
rect 39356 20556 41696 20584
rect 39356 20544 39362 20556
rect 41690 20544 41696 20556
rect 41748 20584 41754 20596
rect 41874 20584 41880 20596
rect 41748 20556 41880 20584
rect 41748 20544 41754 20556
rect 41874 20544 41880 20556
rect 41932 20544 41938 20596
rect 44637 20587 44695 20593
rect 44637 20553 44649 20587
rect 44683 20584 44695 20587
rect 45462 20584 45468 20596
rect 44683 20556 45468 20584
rect 44683 20553 44695 20556
rect 44637 20547 44695 20553
rect 45462 20544 45468 20556
rect 45520 20544 45526 20596
rect 35866 20488 37688 20516
rect 33781 20451 33839 20457
rect 33781 20417 33793 20451
rect 33827 20417 33839 20451
rect 33781 20411 33839 20417
rect 28350 20340 28356 20392
rect 28408 20380 28414 20392
rect 28445 20383 28503 20389
rect 28445 20380 28457 20383
rect 28408 20352 28457 20380
rect 28408 20340 28414 20352
rect 28445 20349 28457 20352
rect 28491 20349 28503 20383
rect 28445 20343 28503 20349
rect 31754 20340 31760 20392
rect 31812 20380 31818 20392
rect 33796 20380 33824 20411
rect 33870 20408 33876 20460
rect 33928 20448 33934 20460
rect 34037 20451 34095 20457
rect 34037 20448 34049 20451
rect 33928 20420 34049 20448
rect 33928 20408 33934 20420
rect 34037 20417 34049 20420
rect 34083 20417 34095 20451
rect 34037 20411 34095 20417
rect 34974 20408 34980 20460
rect 35032 20448 35038 20460
rect 35621 20451 35679 20457
rect 35621 20448 35633 20451
rect 35032 20420 35633 20448
rect 35032 20408 35038 20420
rect 35621 20417 35633 20420
rect 35667 20417 35679 20451
rect 35621 20411 35679 20417
rect 37458 20408 37464 20460
rect 37516 20448 37522 20460
rect 37660 20457 37688 20488
rect 42150 20476 42156 20528
rect 42208 20516 42214 20528
rect 45554 20516 45560 20528
rect 42208 20488 45560 20516
rect 42208 20476 42214 20488
rect 45554 20476 45560 20488
rect 45612 20476 45618 20528
rect 37553 20451 37611 20457
rect 37553 20448 37565 20451
rect 37516 20420 37565 20448
rect 37516 20408 37522 20420
rect 37553 20417 37565 20420
rect 37599 20417 37611 20451
rect 37553 20411 37611 20417
rect 37645 20451 37703 20457
rect 37645 20417 37657 20451
rect 37691 20417 37703 20451
rect 37645 20411 37703 20417
rect 37737 20451 37795 20457
rect 37737 20417 37749 20451
rect 37783 20417 37795 20451
rect 37737 20411 37795 20417
rect 31812 20352 33824 20380
rect 31812 20340 31818 20352
rect 37182 20340 37188 20392
rect 37240 20380 37246 20392
rect 37752 20380 37780 20411
rect 37826 20408 37832 20460
rect 37884 20448 37890 20460
rect 37921 20451 37979 20457
rect 37921 20448 37933 20451
rect 37884 20420 37933 20448
rect 37884 20408 37890 20420
rect 37921 20417 37933 20420
rect 37967 20417 37979 20451
rect 39114 20448 39120 20460
rect 39075 20420 39120 20448
rect 37921 20411 37979 20417
rect 39114 20408 39120 20420
rect 39172 20408 39178 20460
rect 39393 20451 39451 20457
rect 39393 20417 39405 20451
rect 39439 20448 39451 20451
rect 39482 20448 39488 20460
rect 39439 20420 39488 20448
rect 39439 20417 39451 20420
rect 39393 20411 39451 20417
rect 37240 20352 37780 20380
rect 37240 20340 37246 20352
rect 38194 20340 38200 20392
rect 38252 20380 38258 20392
rect 39408 20380 39436 20411
rect 39482 20408 39488 20420
rect 39540 20408 39546 20460
rect 44818 20448 44824 20460
rect 44779 20420 44824 20448
rect 44818 20408 44824 20420
rect 44876 20408 44882 20460
rect 44910 20408 44916 20460
rect 44968 20448 44974 20460
rect 45097 20451 45155 20457
rect 45097 20448 45109 20451
rect 44968 20420 45109 20448
rect 44968 20408 44974 20420
rect 45097 20417 45109 20420
rect 45143 20417 45155 20451
rect 45097 20411 45155 20417
rect 46566 20408 46572 20460
rect 46624 20448 46630 20460
rect 47581 20451 47639 20457
rect 47581 20448 47593 20451
rect 46624 20420 47593 20448
rect 46624 20408 46630 20420
rect 47581 20417 47593 20420
rect 47627 20417 47639 20451
rect 47581 20411 47639 20417
rect 38252 20352 39436 20380
rect 38252 20340 38258 20352
rect 44726 20340 44732 20392
rect 44784 20380 44790 20392
rect 45005 20383 45063 20389
rect 45005 20380 45017 20383
rect 44784 20352 45017 20380
rect 44784 20340 44790 20352
rect 45005 20349 45017 20352
rect 45051 20349 45063 20383
rect 45005 20343 45063 20349
rect 27709 20275 27767 20281
rect 28092 20284 28212 20312
rect 25866 20244 25872 20256
rect 25827 20216 25872 20244
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 27525 20247 27583 20253
rect 27525 20213 27537 20247
rect 27571 20244 27583 20247
rect 28092 20244 28120 20284
rect 35342 20272 35348 20324
rect 35400 20312 35406 20324
rect 38378 20312 38384 20324
rect 35400 20284 38384 20312
rect 35400 20272 35406 20284
rect 38378 20272 38384 20284
rect 38436 20272 38442 20324
rect 28258 20244 28264 20256
rect 27571 20216 28120 20244
rect 28171 20216 28264 20244
rect 27571 20213 27583 20216
rect 27525 20207 27583 20213
rect 28258 20204 28264 20216
rect 28316 20244 28322 20256
rect 30282 20244 30288 20256
rect 28316 20216 30288 20244
rect 28316 20204 28322 20216
rect 30282 20204 30288 20216
rect 30340 20204 30346 20256
rect 33045 20247 33103 20253
rect 33045 20213 33057 20247
rect 33091 20244 33103 20247
rect 33686 20244 33692 20256
rect 33091 20216 33692 20244
rect 33091 20213 33103 20216
rect 33045 20207 33103 20213
rect 33686 20204 33692 20216
rect 33744 20204 33750 20256
rect 34698 20204 34704 20256
rect 34756 20244 34762 20256
rect 35161 20247 35219 20253
rect 35161 20244 35173 20247
rect 34756 20216 35173 20244
rect 34756 20204 34762 20216
rect 35161 20213 35173 20216
rect 35207 20244 35219 20247
rect 35618 20244 35624 20256
rect 35207 20216 35624 20244
rect 35207 20213 35219 20216
rect 35161 20207 35219 20213
rect 35618 20204 35624 20216
rect 35676 20204 35682 20256
rect 36354 20204 36360 20256
rect 36412 20244 36418 20256
rect 38933 20247 38991 20253
rect 38933 20244 38945 20247
rect 36412 20216 38945 20244
rect 36412 20204 36418 20216
rect 38933 20213 38945 20216
rect 38979 20213 38991 20247
rect 38933 20207 38991 20213
rect 39301 20247 39359 20253
rect 39301 20213 39313 20247
rect 39347 20244 39359 20247
rect 41874 20244 41880 20256
rect 39347 20216 41880 20244
rect 39347 20213 39359 20216
rect 39301 20207 39359 20213
rect 41874 20204 41880 20216
rect 41932 20204 41938 20256
rect 46474 20204 46480 20256
rect 46532 20244 46538 20256
rect 47673 20247 47731 20253
rect 47673 20244 47685 20247
rect 46532 20216 47685 20244
rect 46532 20204 46538 20216
rect 47673 20213 47685 20216
rect 47719 20213 47731 20247
rect 47673 20207 47731 20213
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 2590 20040 2596 20052
rect 2551 20012 2596 20040
rect 2590 20000 2596 20012
rect 2648 20000 2654 20052
rect 26237 20043 26295 20049
rect 26237 20009 26249 20043
rect 26283 20040 26295 20043
rect 26326 20040 26332 20052
rect 26283 20012 26332 20040
rect 26283 20009 26295 20012
rect 26237 20003 26295 20009
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 27338 20000 27344 20052
rect 27396 20040 27402 20052
rect 28077 20043 28135 20049
rect 28077 20040 28089 20043
rect 27396 20012 28089 20040
rect 27396 20000 27402 20012
rect 28077 20009 28089 20012
rect 28123 20009 28135 20043
rect 30190 20040 30196 20052
rect 30151 20012 30196 20040
rect 28077 20003 28135 20009
rect 30190 20000 30196 20012
rect 30248 20000 30254 20052
rect 33781 20043 33839 20049
rect 33781 20009 33793 20043
rect 33827 20040 33839 20043
rect 33870 20040 33876 20052
rect 33827 20012 33876 20040
rect 33827 20009 33839 20012
rect 33781 20003 33839 20009
rect 33870 20000 33876 20012
rect 33928 20000 33934 20052
rect 34885 20043 34943 20049
rect 34885 20009 34897 20043
rect 34931 20009 34943 20043
rect 34885 20003 34943 20009
rect 35069 20043 35127 20049
rect 35069 20009 35081 20043
rect 35115 20040 35127 20043
rect 35342 20040 35348 20052
rect 35115 20012 35348 20040
rect 35115 20009 35127 20012
rect 35069 20003 35127 20009
rect 30285 19975 30343 19981
rect 30285 19941 30297 19975
rect 30331 19972 30343 19975
rect 31018 19972 31024 19984
rect 30331 19944 31024 19972
rect 30331 19941 30343 19944
rect 30285 19935 30343 19941
rect 31018 19932 31024 19944
rect 31076 19932 31082 19984
rect 33686 19972 33692 19984
rect 33647 19944 33692 19972
rect 33686 19932 33692 19944
rect 33744 19932 33750 19984
rect 24854 19904 24860 19916
rect 24815 19876 24860 19904
rect 24854 19864 24860 19876
rect 24912 19864 24918 19916
rect 31754 19904 31760 19916
rect 31715 19876 31760 19904
rect 31754 19864 31760 19876
rect 31812 19864 31818 19916
rect 33226 19864 33232 19916
rect 33284 19904 33290 19916
rect 34422 19904 34428 19916
rect 33284 19876 34428 19904
rect 33284 19864 33290 19876
rect 34422 19864 34428 19876
rect 34480 19904 34486 19916
rect 34900 19904 34928 20003
rect 34480 19876 34928 19904
rect 34480 19864 34486 19876
rect 2501 19839 2559 19845
rect 2501 19805 2513 19839
rect 2547 19836 2559 19839
rect 17310 19836 17316 19848
rect 2547 19808 17316 19836
rect 2547 19805 2559 19808
rect 2501 19799 2559 19805
rect 2516 19712 2544 19799
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 24872 19836 24900 19864
rect 26697 19839 26755 19845
rect 26697 19836 26709 19839
rect 24872 19808 26709 19836
rect 26697 19805 26709 19808
rect 26743 19805 26755 19839
rect 26697 19799 26755 19805
rect 30193 19839 30251 19845
rect 30193 19805 30205 19839
rect 30239 19836 30251 19839
rect 30282 19836 30288 19848
rect 30239 19808 30288 19836
rect 30239 19805 30251 19808
rect 30193 19799 30251 19805
rect 30282 19796 30288 19808
rect 30340 19796 30346 19848
rect 30469 19839 30527 19845
rect 30469 19805 30481 19839
rect 30515 19836 30527 19839
rect 31846 19836 31852 19848
rect 30515 19808 31852 19836
rect 30515 19805 30527 19808
rect 30469 19799 30527 19805
rect 31846 19796 31852 19808
rect 31904 19836 31910 19848
rect 32490 19836 32496 19848
rect 31904 19808 32496 19836
rect 31904 19796 31910 19808
rect 32490 19796 32496 19808
rect 32548 19796 32554 19848
rect 33597 19839 33655 19845
rect 33597 19805 33609 19839
rect 33643 19836 33655 19839
rect 35084 19836 35112 20003
rect 35342 20000 35348 20012
rect 35400 20000 35406 20052
rect 37458 20040 37464 20052
rect 37419 20012 37464 20040
rect 37458 20000 37464 20012
rect 37516 20000 37522 20052
rect 40494 20000 40500 20052
rect 40552 20040 40558 20052
rect 41506 20040 41512 20052
rect 40552 20012 41512 20040
rect 40552 20000 40558 20012
rect 41506 20000 41512 20012
rect 41564 20040 41570 20052
rect 41601 20043 41659 20049
rect 41601 20040 41613 20043
rect 41564 20012 41613 20040
rect 41564 20000 41570 20012
rect 41601 20009 41613 20012
rect 41647 20009 41659 20043
rect 41601 20003 41659 20009
rect 45462 20000 45468 20052
rect 45520 20040 45526 20052
rect 45557 20043 45615 20049
rect 45557 20040 45569 20043
rect 45520 20012 45569 20040
rect 45520 20000 45526 20012
rect 45557 20009 45569 20012
rect 45603 20009 45615 20043
rect 45557 20003 45615 20009
rect 35434 19864 35440 19916
rect 35492 19904 35498 19916
rect 36081 19907 36139 19913
rect 36081 19904 36093 19907
rect 35492 19876 36093 19904
rect 35492 19864 35498 19876
rect 36081 19873 36093 19876
rect 36127 19873 36139 19907
rect 36081 19867 36139 19873
rect 36354 19845 36360 19848
rect 36348 19836 36360 19845
rect 33643 19808 35112 19836
rect 36315 19808 36360 19836
rect 33643 19805 33655 19808
rect 33597 19799 33655 19805
rect 36348 19799 36360 19808
rect 36354 19796 36360 19799
rect 36412 19796 36418 19848
rect 37476 19836 37504 20000
rect 38194 19972 38200 19984
rect 38155 19944 38200 19972
rect 38194 19932 38200 19944
rect 38252 19932 38258 19984
rect 39298 19904 39304 19916
rect 38764 19876 39304 19904
rect 38764 19845 38792 19876
rect 39298 19864 39304 19876
rect 39356 19864 39362 19916
rect 42058 19904 42064 19916
rect 41386 19876 42064 19904
rect 38013 19839 38071 19845
rect 38013 19836 38025 19839
rect 37476 19808 38025 19836
rect 38013 19805 38025 19808
rect 38059 19805 38071 19839
rect 38013 19799 38071 19805
rect 38749 19839 38807 19845
rect 38749 19805 38761 19839
rect 38795 19805 38807 19839
rect 38749 19799 38807 19805
rect 38933 19839 38991 19845
rect 38933 19805 38945 19839
rect 38979 19836 38991 19839
rect 39114 19836 39120 19848
rect 38979 19808 39120 19836
rect 38979 19805 38991 19808
rect 38933 19799 38991 19805
rect 39114 19796 39120 19808
rect 39172 19836 39178 19848
rect 39666 19836 39672 19848
rect 39172 19808 39672 19836
rect 39172 19796 39178 19808
rect 39666 19796 39672 19808
rect 39724 19796 39730 19848
rect 40218 19836 40224 19848
rect 40179 19808 40224 19836
rect 40218 19796 40224 19808
rect 40276 19836 40282 19848
rect 41386 19836 41414 19876
rect 42058 19864 42064 19876
rect 42116 19864 42122 19916
rect 43254 19864 43260 19916
rect 43312 19904 43318 19916
rect 44450 19904 44456 19916
rect 43312 19876 44456 19904
rect 43312 19864 43318 19876
rect 44450 19864 44456 19876
rect 44508 19904 44514 19916
rect 46474 19904 46480 19916
rect 44508 19876 45324 19904
rect 46435 19876 46480 19904
rect 44508 19864 44514 19876
rect 45296 19848 45324 19876
rect 46474 19864 46480 19876
rect 46532 19864 46538 19916
rect 48130 19904 48136 19916
rect 48091 19876 48136 19904
rect 48130 19864 48136 19876
rect 48188 19864 48194 19916
rect 40276 19808 41414 19836
rect 44269 19839 44327 19845
rect 40276 19796 40282 19808
rect 44269 19805 44281 19839
rect 44315 19836 44327 19839
rect 44818 19836 44824 19848
rect 44315 19808 44824 19836
rect 44315 19805 44327 19808
rect 44269 19799 44327 19805
rect 44818 19796 44824 19808
rect 44876 19796 44882 19848
rect 45278 19796 45284 19848
rect 45336 19836 45342 19848
rect 45465 19839 45523 19845
rect 45465 19836 45477 19839
rect 45336 19808 45477 19836
rect 45336 19796 45342 19808
rect 45465 19805 45477 19808
rect 45511 19805 45523 19839
rect 45465 19799 45523 19805
rect 46293 19839 46351 19845
rect 46293 19805 46305 19839
rect 46339 19805 46351 19839
rect 46293 19799 46351 19805
rect 25124 19771 25182 19777
rect 25124 19737 25136 19771
rect 25170 19768 25182 19771
rect 25866 19768 25872 19780
rect 25170 19740 25872 19768
rect 25170 19737 25182 19740
rect 25124 19731 25182 19737
rect 25866 19728 25872 19740
rect 25924 19728 25930 19780
rect 26964 19771 27022 19777
rect 26964 19737 26976 19771
rect 27010 19768 27022 19771
rect 27154 19768 27160 19780
rect 27010 19740 27160 19768
rect 27010 19737 27022 19740
rect 26964 19731 27022 19737
rect 27154 19728 27160 19740
rect 27212 19728 27218 19780
rect 32024 19771 32082 19777
rect 32024 19737 32036 19771
rect 32070 19768 32082 19771
rect 32398 19768 32404 19780
rect 32070 19740 32404 19768
rect 32070 19737 32082 19740
rect 32024 19731 32082 19737
rect 32398 19728 32404 19740
rect 32456 19728 32462 19780
rect 32508 19768 32536 19796
rect 33873 19771 33931 19777
rect 33873 19768 33885 19771
rect 32508 19740 33885 19768
rect 33873 19737 33885 19740
rect 33919 19737 33931 19771
rect 34698 19768 34704 19780
rect 34659 19740 34704 19768
rect 33873 19731 33931 19737
rect 34698 19728 34704 19740
rect 34756 19728 34762 19780
rect 37182 19728 37188 19780
rect 37240 19768 37246 19780
rect 37240 19740 40264 19768
rect 37240 19728 37246 19740
rect 2498 19660 2504 19712
rect 2556 19660 2562 19712
rect 32306 19660 32312 19712
rect 32364 19700 32370 19712
rect 33137 19703 33195 19709
rect 33137 19700 33149 19703
rect 32364 19672 33149 19700
rect 32364 19660 32370 19672
rect 33137 19669 33149 19672
rect 33183 19700 33195 19703
rect 33410 19700 33416 19712
rect 33183 19672 33416 19700
rect 33183 19669 33195 19672
rect 33137 19663 33195 19669
rect 33410 19660 33416 19672
rect 33468 19700 33474 19712
rect 34790 19700 34796 19712
rect 33468 19672 34796 19700
rect 33468 19660 33474 19672
rect 34790 19660 34796 19672
rect 34848 19700 34854 19712
rect 34901 19703 34959 19709
rect 34901 19700 34913 19703
rect 34848 19672 34913 19700
rect 34848 19660 34854 19672
rect 34901 19669 34913 19672
rect 34947 19669 34959 19703
rect 38838 19700 38844 19712
rect 38799 19672 38844 19700
rect 34901 19663 34959 19669
rect 38838 19660 38844 19672
rect 38896 19660 38902 19712
rect 40236 19700 40264 19740
rect 40310 19728 40316 19780
rect 40368 19768 40374 19780
rect 42334 19777 42340 19780
rect 40466 19771 40524 19777
rect 40466 19768 40478 19771
rect 40368 19740 40478 19768
rect 40368 19728 40374 19740
rect 40466 19737 40478 19740
rect 40512 19737 40524 19771
rect 40466 19731 40524 19737
rect 42328 19731 42340 19777
rect 42392 19768 42398 19780
rect 45186 19768 45192 19780
rect 42392 19740 42428 19768
rect 42536 19740 45192 19768
rect 42334 19728 42340 19731
rect 42392 19728 42398 19740
rect 40862 19700 40868 19712
rect 40236 19672 40868 19700
rect 40862 19660 40868 19672
rect 40920 19700 40926 19712
rect 42536 19700 42564 19740
rect 45186 19728 45192 19740
rect 45244 19728 45250 19780
rect 46308 19768 46336 19799
rect 47762 19768 47768 19780
rect 46308 19740 47768 19768
rect 47762 19728 47768 19740
rect 47820 19728 47826 19780
rect 40920 19672 42564 19700
rect 40920 19660 40926 19672
rect 42610 19660 42616 19712
rect 42668 19700 42674 19712
rect 43441 19703 43499 19709
rect 43441 19700 43453 19703
rect 42668 19672 43453 19700
rect 42668 19660 42674 19672
rect 43441 19669 43453 19672
rect 43487 19700 43499 19703
rect 43622 19700 43628 19712
rect 43487 19672 43628 19700
rect 43487 19669 43499 19672
rect 43441 19663 43499 19669
rect 43622 19660 43628 19672
rect 43680 19660 43686 19712
rect 44358 19700 44364 19712
rect 44319 19672 44364 19700
rect 44358 19660 44364 19672
rect 44416 19660 44422 19712
rect 45204 19700 45232 19728
rect 46290 19700 46296 19712
rect 45204 19672 46296 19700
rect 46290 19660 46296 19672
rect 46348 19660 46354 19712
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 27154 19496 27160 19508
rect 27115 19468 27160 19496
rect 27154 19456 27160 19468
rect 27212 19456 27218 19508
rect 32398 19496 32404 19508
rect 32359 19468 32404 19496
rect 32398 19456 32404 19468
rect 32456 19456 32462 19508
rect 34422 19496 34428 19508
rect 34383 19468 34428 19496
rect 34422 19456 34428 19468
rect 34480 19456 34486 19508
rect 37826 19456 37832 19508
rect 37884 19496 37890 19508
rect 39209 19499 39267 19505
rect 39209 19496 39221 19499
rect 37884 19468 39221 19496
rect 37884 19456 37890 19468
rect 39209 19465 39221 19468
rect 39255 19465 39267 19499
rect 39209 19459 39267 19465
rect 44545 19499 44603 19505
rect 44545 19465 44557 19499
rect 44591 19496 44603 19499
rect 44591 19468 45937 19496
rect 44591 19465 44603 19468
rect 44545 19459 44603 19465
rect 31754 19388 31760 19440
rect 31812 19428 31818 19440
rect 33318 19437 33324 19440
rect 33312 19428 33324 19437
rect 31812 19400 33088 19428
rect 33279 19400 33324 19428
rect 31812 19388 31818 19400
rect 27062 19360 27068 19372
rect 27023 19332 27068 19360
rect 27062 19320 27068 19332
rect 27120 19320 27126 19372
rect 27246 19360 27252 19372
rect 27207 19332 27252 19360
rect 27246 19320 27252 19332
rect 27304 19320 27310 19372
rect 32306 19360 32312 19372
rect 32267 19332 32312 19360
rect 32306 19320 32312 19332
rect 32364 19320 32370 19372
rect 32490 19360 32496 19372
rect 32451 19332 32496 19360
rect 32490 19320 32496 19332
rect 32548 19320 32554 19372
rect 33060 19369 33088 19400
rect 33312 19391 33324 19400
rect 33318 19388 33324 19391
rect 33376 19388 33382 19440
rect 33778 19388 33784 19440
rect 33836 19428 33842 19440
rect 37182 19428 37188 19440
rect 33836 19400 37188 19428
rect 33836 19388 33842 19400
rect 37182 19388 37188 19400
rect 37240 19388 37246 19440
rect 40218 19428 40224 19440
rect 37292 19400 40224 19428
rect 37292 19369 37320 19400
rect 40218 19388 40224 19400
rect 40276 19388 40282 19440
rect 40770 19428 40776 19440
rect 40696 19400 40776 19428
rect 33045 19363 33103 19369
rect 33045 19329 33057 19363
rect 33091 19329 33103 19363
rect 33045 19323 33103 19329
rect 37277 19363 37335 19369
rect 37277 19329 37289 19363
rect 37323 19329 37335 19363
rect 37277 19323 37335 19329
rect 37544 19363 37602 19369
rect 37544 19329 37556 19363
rect 37590 19360 37602 19363
rect 38746 19360 38752 19372
rect 37590 19332 38752 19360
rect 37590 19329 37602 19332
rect 37544 19323 37602 19329
rect 38746 19320 38752 19332
rect 38804 19320 38810 19372
rect 39114 19360 39120 19372
rect 39075 19332 39120 19360
rect 39114 19320 39120 19332
rect 39172 19320 39178 19372
rect 40310 19360 40316 19372
rect 40236 19332 40316 19360
rect 38657 19227 38715 19233
rect 38657 19193 38669 19227
rect 38703 19224 38715 19227
rect 39132 19224 39160 19320
rect 40236 19301 40264 19332
rect 40310 19320 40316 19332
rect 40368 19320 40374 19372
rect 40402 19320 40408 19372
rect 40460 19369 40466 19372
rect 40696 19369 40724 19400
rect 40770 19388 40776 19400
rect 40828 19388 40834 19440
rect 41690 19428 41696 19440
rect 41603 19400 41696 19428
rect 41690 19388 41696 19400
rect 41748 19428 41754 19440
rect 45909 19437 45937 19468
rect 46014 19456 46020 19508
rect 46072 19496 46078 19508
rect 47029 19499 47087 19505
rect 47029 19496 47041 19499
rect 46072 19468 47041 19496
rect 46072 19456 46078 19468
rect 47029 19465 47041 19468
rect 47075 19465 47087 19499
rect 47029 19459 47087 19465
rect 45894 19431 45952 19437
rect 41748 19400 43576 19428
rect 41748 19388 41754 19400
rect 40460 19363 40509 19369
rect 40460 19329 40463 19363
rect 40497 19329 40509 19363
rect 40460 19323 40509 19329
rect 40586 19363 40644 19369
rect 40586 19329 40598 19363
rect 40632 19329 40644 19363
rect 40586 19323 40644 19329
rect 40681 19363 40739 19369
rect 40681 19329 40693 19363
rect 40727 19329 40739 19363
rect 40681 19323 40739 19329
rect 40460 19320 40466 19323
rect 40221 19295 40279 19301
rect 40221 19261 40233 19295
rect 40267 19261 40279 19295
rect 40221 19255 40279 19261
rect 38703 19196 39160 19224
rect 40604 19224 40632 19323
rect 40862 19320 40868 19372
rect 40920 19360 40926 19372
rect 42444 19369 42472 19400
rect 42429 19363 42487 19369
rect 40920 19332 40965 19360
rect 40920 19320 40926 19332
rect 42429 19329 42441 19363
rect 42475 19329 42487 19363
rect 42610 19360 42616 19372
rect 42571 19332 42616 19360
rect 42429 19323 42487 19329
rect 42610 19320 42616 19332
rect 42668 19320 42674 19372
rect 43254 19360 43260 19372
rect 43215 19332 43260 19360
rect 43254 19320 43260 19332
rect 43312 19320 43318 19372
rect 43548 19369 43576 19400
rect 45894 19397 45906 19431
rect 45940 19397 45952 19431
rect 45894 19391 45952 19397
rect 43533 19363 43591 19369
rect 43533 19329 43545 19363
rect 43579 19329 43591 19363
rect 43533 19323 43591 19329
rect 44634 19320 44640 19372
rect 44692 19360 44698 19372
rect 44775 19363 44833 19369
rect 44775 19360 44787 19363
rect 44692 19332 44787 19360
rect 44692 19320 44698 19332
rect 44775 19329 44787 19332
rect 44821 19329 44833 19363
rect 44775 19323 44833 19329
rect 44910 19363 44968 19369
rect 44910 19329 44922 19363
rect 44956 19329 44968 19363
rect 44910 19323 44968 19329
rect 44928 19292 44956 19323
rect 45002 19320 45008 19372
rect 45060 19369 45066 19372
rect 45060 19360 45068 19369
rect 45060 19332 45105 19360
rect 45060 19323 45068 19332
rect 45060 19320 45066 19323
rect 45186 19320 45192 19372
rect 45244 19360 45250 19372
rect 45649 19363 45707 19369
rect 45244 19332 45289 19360
rect 45244 19320 45250 19332
rect 45649 19329 45661 19363
rect 45695 19360 45707 19363
rect 46750 19360 46756 19372
rect 45695 19332 46756 19360
rect 45695 19329 45707 19332
rect 45649 19323 45707 19329
rect 46750 19320 46756 19332
rect 46808 19320 46814 19372
rect 47762 19292 47768 19304
rect 44928 19264 45048 19292
rect 47723 19264 47768 19292
rect 41874 19224 41880 19236
rect 40604 19196 41880 19224
rect 38703 19193 38715 19196
rect 38657 19187 38715 19193
rect 41874 19184 41880 19196
rect 41932 19224 41938 19236
rect 41932 19196 43116 19224
rect 41932 19184 41938 19196
rect 42058 19116 42064 19168
rect 42116 19156 42122 19168
rect 42429 19159 42487 19165
rect 42429 19156 42441 19159
rect 42116 19128 42441 19156
rect 42116 19116 42122 19128
rect 42429 19125 42441 19128
rect 42475 19125 42487 19159
rect 43088 19156 43116 19196
rect 45020 19156 45048 19264
rect 47762 19252 47768 19264
rect 47820 19252 47826 19304
rect 45922 19156 45928 19168
rect 43088 19128 45928 19156
rect 42429 19119 42487 19125
rect 45922 19116 45928 19128
rect 45980 19116 45986 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 38657 18955 38715 18961
rect 38657 18921 38669 18955
rect 38703 18952 38715 18955
rect 38838 18952 38844 18964
rect 38703 18924 38844 18952
rect 38703 18921 38715 18924
rect 38657 18915 38715 18921
rect 38838 18912 38844 18924
rect 38896 18912 38902 18964
rect 40497 18955 40555 18961
rect 40497 18921 40509 18955
rect 40543 18952 40555 18955
rect 40770 18952 40776 18964
rect 40543 18924 40776 18952
rect 40543 18921 40555 18924
rect 40497 18915 40555 18921
rect 40770 18912 40776 18924
rect 40828 18912 40834 18964
rect 42058 18952 42064 18964
rect 42019 18924 42064 18952
rect 42058 18912 42064 18924
rect 42116 18912 42122 18964
rect 42245 18955 42303 18961
rect 42245 18921 42257 18955
rect 42291 18952 42303 18955
rect 42334 18952 42340 18964
rect 42291 18924 42340 18952
rect 42291 18921 42303 18924
rect 42245 18915 42303 18921
rect 42334 18912 42340 18924
rect 42392 18912 42398 18964
rect 43530 18952 43536 18964
rect 42904 18924 43536 18952
rect 38746 18884 38752 18896
rect 38707 18856 38752 18884
rect 38746 18844 38752 18856
rect 38804 18844 38810 18896
rect 40034 18844 40040 18896
rect 40092 18884 40098 18896
rect 42904 18884 42932 18924
rect 43530 18912 43536 18924
rect 43588 18952 43594 18964
rect 44634 18952 44640 18964
rect 43588 18924 44640 18952
rect 43588 18912 43594 18924
rect 44634 18912 44640 18924
rect 44692 18952 44698 18964
rect 45235 18955 45293 18961
rect 45235 18952 45247 18955
rect 44692 18924 45247 18952
rect 44692 18912 44698 18924
rect 45235 18921 45247 18924
rect 45281 18921 45293 18955
rect 45235 18915 45293 18921
rect 44358 18884 44364 18896
rect 40092 18856 42932 18884
rect 43364 18856 44364 18884
rect 40092 18844 40098 18856
rect 41598 18816 41604 18828
rect 38764 18788 41604 18816
rect 2130 18708 2136 18760
rect 2188 18748 2194 18760
rect 2317 18751 2375 18757
rect 2317 18748 2329 18751
rect 2188 18720 2329 18748
rect 2188 18708 2194 18720
rect 2317 18717 2329 18720
rect 2363 18717 2375 18751
rect 2317 18711 2375 18717
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18748 2835 18751
rect 2866 18748 2872 18760
rect 2823 18720 2872 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 38764 18757 38792 18788
rect 41598 18776 41604 18788
rect 41656 18816 41662 18828
rect 42153 18819 42211 18825
rect 42153 18816 42165 18819
rect 41656 18788 42165 18816
rect 41656 18776 41662 18788
rect 42153 18785 42165 18788
rect 42199 18785 42211 18819
rect 42153 18779 42211 18785
rect 38749 18751 38807 18757
rect 38749 18717 38761 18751
rect 38795 18717 38807 18751
rect 40402 18748 40408 18760
rect 40363 18720 40408 18748
rect 38749 18711 38807 18717
rect 40402 18708 40408 18720
rect 40460 18708 40466 18760
rect 40589 18751 40647 18757
rect 40589 18717 40601 18751
rect 40635 18748 40647 18751
rect 41969 18751 42027 18757
rect 41969 18748 41981 18751
rect 40635 18720 41981 18748
rect 40635 18717 40647 18720
rect 40589 18711 40647 18717
rect 41969 18717 41981 18720
rect 42015 18748 42027 18751
rect 42058 18748 42064 18760
rect 42015 18720 42064 18748
rect 42015 18717 42027 18720
rect 41969 18711 42027 18717
rect 38381 18683 38439 18689
rect 38381 18649 38393 18683
rect 38427 18680 38439 18683
rect 39206 18680 39212 18692
rect 38427 18652 39212 18680
rect 38427 18649 38439 18652
rect 38381 18643 38439 18649
rect 39206 18640 39212 18652
rect 39264 18640 39270 18692
rect 2314 18572 2320 18624
rect 2372 18612 2378 18624
rect 2869 18615 2927 18621
rect 2869 18612 2881 18615
rect 2372 18584 2881 18612
rect 2372 18572 2378 18584
rect 2869 18581 2881 18584
rect 2915 18581 2927 18615
rect 2869 18575 2927 18581
rect 38473 18615 38531 18621
rect 38473 18581 38485 18615
rect 38519 18612 38531 18615
rect 40604 18612 40632 18711
rect 42058 18708 42064 18720
rect 42116 18708 42122 18760
rect 42610 18708 42616 18760
rect 42668 18748 42674 18760
rect 43364 18757 43392 18856
rect 44358 18844 44364 18856
rect 44416 18884 44422 18896
rect 45462 18884 45468 18896
rect 44416 18856 45468 18884
rect 44416 18844 44422 18856
rect 45462 18844 45468 18856
rect 45520 18844 45526 18896
rect 43622 18816 43628 18828
rect 43583 18788 43628 18816
rect 43622 18776 43628 18788
rect 43680 18776 43686 18828
rect 45005 18819 45063 18825
rect 45005 18785 45017 18819
rect 45051 18816 45063 18819
rect 46014 18816 46020 18828
rect 45051 18788 46020 18816
rect 45051 18785 45063 18788
rect 45005 18779 45063 18785
rect 46014 18776 46020 18788
rect 46072 18776 46078 18828
rect 48130 18816 48136 18828
rect 48091 18788 48136 18816
rect 48130 18776 48136 18788
rect 48188 18776 48194 18828
rect 43349 18751 43407 18757
rect 43349 18748 43361 18751
rect 42668 18720 43361 18748
rect 42668 18708 42674 18720
rect 43349 18717 43361 18720
rect 43395 18717 43407 18751
rect 44266 18748 44272 18760
rect 44227 18720 44272 18748
rect 43349 18711 43407 18717
rect 44266 18708 44272 18720
rect 44324 18708 44330 18760
rect 46290 18748 46296 18760
rect 46251 18720 46296 18748
rect 46290 18708 46296 18720
rect 46348 18708 46354 18760
rect 41785 18683 41843 18689
rect 41785 18649 41797 18683
rect 41831 18680 41843 18683
rect 43070 18680 43076 18692
rect 41831 18652 43076 18680
rect 41831 18649 41843 18652
rect 41785 18643 41843 18649
rect 43070 18640 43076 18652
rect 43128 18640 43134 18692
rect 44082 18680 44088 18692
rect 44043 18652 44088 18680
rect 44082 18640 44088 18652
rect 44140 18640 44146 18692
rect 46477 18683 46535 18689
rect 46477 18649 46489 18683
rect 46523 18680 46535 18683
rect 46934 18680 46940 18692
rect 46523 18652 46940 18680
rect 46523 18649 46535 18652
rect 46477 18643 46535 18649
rect 46934 18640 46940 18652
rect 46992 18640 46998 18692
rect 43162 18612 43168 18624
rect 38519 18584 40632 18612
rect 43123 18584 43168 18612
rect 38519 18581 38531 18584
rect 38473 18575 38531 18581
rect 43162 18572 43168 18584
rect 43220 18572 43226 18624
rect 44453 18615 44511 18621
rect 44453 18581 44465 18615
rect 44499 18612 44511 18615
rect 44726 18612 44732 18624
rect 44499 18584 44732 18612
rect 44499 18581 44511 18584
rect 44453 18575 44511 18581
rect 44726 18572 44732 18584
rect 44784 18572 44790 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 44361 18411 44419 18417
rect 44361 18377 44373 18411
rect 44407 18408 44419 18411
rect 44450 18408 44456 18420
rect 44407 18380 44456 18408
rect 44407 18377 44419 18380
rect 44361 18371 44419 18377
rect 44450 18368 44456 18380
rect 44508 18368 44514 18420
rect 45002 18408 45008 18420
rect 44963 18380 45008 18408
rect 45002 18368 45008 18380
rect 45060 18368 45066 18420
rect 46934 18408 46940 18420
rect 46895 18380 46940 18408
rect 46934 18368 46940 18380
rect 46992 18368 46998 18420
rect 2314 18340 2320 18352
rect 2275 18312 2320 18340
rect 2314 18300 2320 18312
rect 2372 18300 2378 18352
rect 42521 18343 42579 18349
rect 42521 18309 42533 18343
rect 42567 18340 42579 18343
rect 42610 18340 42616 18352
rect 42567 18312 42616 18340
rect 42567 18309 42579 18312
rect 42521 18303 42579 18309
rect 42610 18300 42616 18312
rect 42668 18300 42674 18352
rect 42705 18343 42763 18349
rect 42705 18309 42717 18343
rect 42751 18340 42763 18343
rect 42978 18340 42984 18352
rect 42751 18312 42984 18340
rect 42751 18309 42763 18312
rect 42705 18303 42763 18309
rect 42978 18300 42984 18312
rect 43036 18300 43042 18352
rect 43165 18343 43223 18349
rect 43165 18309 43177 18343
rect 43211 18340 43223 18343
rect 44174 18340 44180 18352
rect 43211 18312 44180 18340
rect 43211 18309 43223 18312
rect 43165 18303 43223 18309
rect 44174 18300 44180 18312
rect 44232 18340 44238 18352
rect 44232 18312 44864 18340
rect 44232 18300 44238 18312
rect 2130 18272 2136 18284
rect 2091 18244 2136 18272
rect 2130 18232 2136 18244
rect 2188 18232 2194 18284
rect 2774 18204 2780 18216
rect 2735 18176 2780 18204
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18204 13047 18207
rect 13449 18207 13507 18213
rect 13449 18204 13461 18207
rect 13035 18176 13461 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 13449 18173 13461 18176
rect 13495 18173 13507 18207
rect 13630 18204 13636 18216
rect 13591 18176 13636 18204
rect 13449 18167 13507 18173
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 15102 18204 15108 18216
rect 15063 18176 15108 18204
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 42426 18164 42432 18216
rect 42484 18204 42490 18216
rect 42996 18204 43024 18300
rect 43530 18272 43536 18284
rect 43491 18244 43536 18272
rect 43530 18232 43536 18244
rect 43588 18232 43594 18284
rect 44726 18272 44732 18284
rect 44687 18244 44732 18272
rect 44726 18232 44732 18244
rect 44784 18232 44790 18284
rect 44836 18281 44864 18312
rect 46290 18300 46296 18352
rect 46348 18340 46354 18352
rect 46348 18312 47808 18340
rect 46348 18300 46354 18312
rect 44821 18275 44879 18281
rect 44821 18241 44833 18275
rect 44867 18241 44879 18275
rect 44821 18235 44879 18241
rect 45649 18275 45707 18281
rect 45649 18241 45661 18275
rect 45695 18272 45707 18275
rect 46014 18272 46020 18284
rect 45695 18244 46020 18272
rect 45695 18241 45707 18244
rect 45649 18235 45707 18241
rect 46014 18232 46020 18244
rect 46072 18232 46078 18284
rect 47780 18281 47808 18312
rect 46845 18275 46903 18281
rect 46845 18241 46857 18275
rect 46891 18241 46903 18275
rect 46845 18235 46903 18241
rect 47765 18275 47823 18281
rect 47765 18241 47777 18275
rect 47811 18241 47823 18275
rect 47765 18235 47823 18241
rect 43625 18207 43683 18213
rect 43625 18204 43637 18207
rect 42484 18176 43637 18204
rect 42484 18164 42490 18176
rect 43625 18173 43637 18176
rect 43671 18173 43683 18207
rect 43625 18167 43683 18173
rect 45462 18164 45468 18216
rect 45520 18204 45526 18216
rect 45557 18207 45615 18213
rect 45557 18204 45569 18207
rect 45520 18176 45569 18204
rect 45520 18164 45526 18176
rect 45557 18173 45569 18176
rect 45603 18173 45615 18207
rect 46860 18204 46888 18235
rect 47854 18204 47860 18216
rect 46860 18176 47860 18204
rect 45557 18167 45615 18173
rect 47854 18164 47860 18176
rect 47912 18164 47918 18216
rect 44082 18096 44088 18148
rect 44140 18136 44146 18148
rect 46017 18139 46075 18145
rect 46017 18136 46029 18139
rect 44140 18108 46029 18136
rect 44140 18096 44146 18108
rect 46017 18105 46029 18108
rect 46063 18105 46075 18139
rect 46017 18099 46075 18105
rect 42886 18028 42892 18080
rect 42944 18068 42950 18080
rect 43809 18071 43867 18077
rect 43809 18068 43821 18071
rect 42944 18040 43821 18068
rect 42944 18028 42950 18040
rect 43809 18037 43821 18040
rect 43855 18037 43867 18071
rect 43809 18031 43867 18037
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 13173 17867 13231 17873
rect 13173 17833 13185 17867
rect 13219 17864 13231 17867
rect 13630 17864 13636 17876
rect 13219 17836 13636 17864
rect 13219 17833 13231 17836
rect 13173 17827 13231 17833
rect 13630 17824 13636 17836
rect 13688 17824 13694 17876
rect 15102 17824 15108 17876
rect 15160 17864 15166 17876
rect 45554 17864 45560 17876
rect 15160 17836 45560 17864
rect 15160 17824 15166 17836
rect 45554 17824 45560 17836
rect 45612 17824 45618 17876
rect 38197 17799 38255 17805
rect 38197 17765 38209 17799
rect 38243 17796 38255 17799
rect 39206 17796 39212 17808
rect 38243 17768 38792 17796
rect 39167 17768 39212 17796
rect 38243 17765 38255 17768
rect 38197 17759 38255 17765
rect 38764 17737 38792 17768
rect 39206 17756 39212 17768
rect 39264 17756 39270 17808
rect 42426 17796 42432 17808
rect 40420 17768 42432 17796
rect 37921 17731 37979 17737
rect 37921 17697 37933 17731
rect 37967 17697 37979 17731
rect 37921 17691 37979 17697
rect 38749 17731 38807 17737
rect 38749 17697 38761 17731
rect 38795 17697 38807 17731
rect 38749 17691 38807 17697
rect 2130 17620 2136 17672
rect 2188 17660 2194 17672
rect 2317 17663 2375 17669
rect 2317 17660 2329 17663
rect 2188 17632 2329 17660
rect 2188 17620 2194 17632
rect 2317 17629 2329 17632
rect 2363 17629 2375 17663
rect 2317 17623 2375 17629
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 13078 17660 13084 17672
rect 12584 17632 13084 17660
rect 12584 17620 12590 17632
rect 13078 17620 13084 17632
rect 13136 17620 13142 17672
rect 37826 17660 37832 17672
rect 37787 17632 37832 17660
rect 37826 17620 37832 17632
rect 37884 17620 37890 17672
rect 37936 17592 37964 17691
rect 38841 17663 38899 17669
rect 38841 17629 38853 17663
rect 38887 17660 38899 17663
rect 39850 17660 39856 17672
rect 38887 17632 39856 17660
rect 38887 17629 38899 17632
rect 38841 17623 38899 17629
rect 39850 17620 39856 17632
rect 39908 17620 39914 17672
rect 40420 17669 40448 17768
rect 42426 17756 42432 17768
rect 42484 17756 42490 17808
rect 42702 17796 42708 17808
rect 42536 17768 42708 17796
rect 40494 17688 40500 17740
rect 40552 17728 40558 17740
rect 41049 17731 41107 17737
rect 41049 17728 41061 17731
rect 40552 17700 41061 17728
rect 40552 17688 40558 17700
rect 40604 17669 40632 17700
rect 41049 17697 41061 17700
rect 41095 17697 41107 17731
rect 41049 17691 41107 17697
rect 40405 17663 40463 17669
rect 40405 17629 40417 17663
rect 40451 17629 40463 17663
rect 40405 17623 40463 17629
rect 40589 17663 40647 17669
rect 40589 17629 40601 17663
rect 40635 17660 40647 17663
rect 41233 17663 41291 17669
rect 40635 17632 40669 17660
rect 40635 17629 40647 17632
rect 40589 17623 40647 17629
rect 41233 17629 41245 17663
rect 41279 17660 41291 17663
rect 42536 17660 42564 17768
rect 42702 17756 42708 17768
rect 42760 17756 42766 17808
rect 43070 17796 43076 17808
rect 43031 17768 43076 17796
rect 43070 17756 43076 17768
rect 43128 17756 43134 17808
rect 42613 17731 42671 17737
rect 42613 17697 42625 17731
rect 42659 17728 42671 17731
rect 42886 17728 42892 17740
rect 42659 17700 42892 17728
rect 42659 17697 42671 17700
rect 42613 17691 42671 17697
rect 42886 17688 42892 17700
rect 42944 17688 42950 17740
rect 43162 17688 43168 17740
rect 43220 17728 43226 17740
rect 43993 17731 44051 17737
rect 43993 17728 44005 17731
rect 43220 17700 44005 17728
rect 43220 17688 43226 17700
rect 43993 17697 44005 17700
rect 44039 17697 44051 17731
rect 43993 17691 44051 17697
rect 41279 17632 42564 17660
rect 42705 17663 42763 17669
rect 41279 17629 41291 17632
rect 41233 17623 41291 17629
rect 42705 17629 42717 17663
rect 42751 17660 42763 17663
rect 42978 17660 42984 17672
rect 42751 17632 42984 17660
rect 42751 17629 42763 17632
rect 42705 17623 42763 17629
rect 40420 17592 40448 17623
rect 42978 17620 42984 17632
rect 43036 17660 43042 17672
rect 43717 17663 43775 17669
rect 43717 17660 43729 17663
rect 43036 17632 43729 17660
rect 43036 17620 43042 17632
rect 43717 17629 43729 17632
rect 43763 17629 43775 17663
rect 43717 17623 43775 17629
rect 43809 17663 43867 17669
rect 43809 17629 43821 17663
rect 43855 17629 43867 17663
rect 43809 17623 43867 17629
rect 43901 17663 43959 17669
rect 43901 17629 43913 17663
rect 43947 17660 43959 17663
rect 44266 17660 44272 17672
rect 43947 17632 44272 17660
rect 43947 17629 43959 17632
rect 43901 17623 43959 17629
rect 37936 17564 40448 17592
rect 40954 17552 40960 17604
rect 41012 17592 41018 17604
rect 41417 17595 41475 17601
rect 41417 17592 41429 17595
rect 41012 17564 41429 17592
rect 41012 17552 41018 17564
rect 41417 17561 41429 17564
rect 41463 17561 41475 17595
rect 43824 17592 43852 17623
rect 44266 17620 44272 17632
rect 44324 17620 44330 17672
rect 44082 17592 44088 17604
rect 41417 17555 41475 17561
rect 42444 17564 43576 17592
rect 43824 17564 44088 17592
rect 40497 17527 40555 17533
rect 40497 17493 40509 17527
rect 40543 17524 40555 17527
rect 41138 17524 41144 17536
rect 40543 17496 41144 17524
rect 40543 17493 40555 17496
rect 40497 17487 40555 17493
rect 41138 17484 41144 17496
rect 41196 17484 41202 17536
rect 41230 17484 41236 17536
rect 41288 17524 41294 17536
rect 42444 17524 42472 17564
rect 43548 17533 43576 17564
rect 44082 17552 44088 17564
rect 44140 17552 44146 17604
rect 41288 17496 42472 17524
rect 43533 17527 43591 17533
rect 41288 17484 41294 17496
rect 43533 17493 43545 17527
rect 43579 17493 43591 17527
rect 43533 17487 43591 17493
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 40402 17280 40408 17332
rect 40460 17320 40466 17332
rect 40497 17323 40555 17329
rect 40497 17320 40509 17323
rect 40460 17292 40509 17320
rect 40460 17280 40466 17292
rect 40497 17289 40509 17292
rect 40543 17289 40555 17323
rect 44174 17320 44180 17332
rect 44135 17292 44180 17320
rect 40497 17283 40555 17289
rect 44174 17280 44180 17292
rect 44232 17280 44238 17332
rect 2130 17184 2136 17196
rect 2091 17156 2136 17184
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 40129 17187 40187 17193
rect 40129 17153 40141 17187
rect 40175 17153 40187 17187
rect 40954 17184 40960 17196
rect 40915 17156 40960 17184
rect 40129 17147 40187 17153
rect 2314 17116 2320 17128
rect 2275 17088 2320 17116
rect 2314 17076 2320 17088
rect 2372 17076 2378 17128
rect 2774 17116 2780 17128
rect 2735 17088 2780 17116
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 40037 17119 40095 17125
rect 40037 17085 40049 17119
rect 40083 17085 40095 17119
rect 40144 17116 40172 17147
rect 40954 17144 40960 17156
rect 41012 17144 41018 17196
rect 41138 17184 41144 17196
rect 41099 17156 41144 17184
rect 41138 17144 41144 17156
rect 41196 17144 41202 17196
rect 42613 17187 42671 17193
rect 42613 17153 42625 17187
rect 42659 17184 42671 17187
rect 43622 17184 43628 17196
rect 42659 17156 43628 17184
rect 42659 17153 42671 17156
rect 42613 17147 42671 17153
rect 43622 17144 43628 17156
rect 43680 17144 43686 17196
rect 44082 17184 44088 17196
rect 44043 17156 44088 17184
rect 44082 17144 44088 17156
rect 44140 17144 44146 17196
rect 44266 17184 44272 17196
rect 44227 17156 44272 17184
rect 44266 17144 44272 17156
rect 44324 17144 44330 17196
rect 46845 17187 46903 17193
rect 46845 17153 46857 17187
rect 46891 17184 46903 17187
rect 47394 17184 47400 17196
rect 46891 17156 47400 17184
rect 46891 17153 46903 17156
rect 46845 17147 46903 17153
rect 47394 17144 47400 17156
rect 47452 17144 47458 17196
rect 40218 17116 40224 17128
rect 40144 17088 40224 17116
rect 40037 17079 40095 17085
rect 40052 17048 40080 17079
rect 40218 17076 40224 17088
rect 40276 17116 40282 17128
rect 41049 17119 41107 17125
rect 41049 17116 41061 17119
rect 40276 17088 41061 17116
rect 40276 17076 40282 17088
rect 41049 17085 41061 17088
rect 41095 17085 41107 17119
rect 42702 17116 42708 17128
rect 42663 17088 42708 17116
rect 41049 17079 41107 17085
rect 42702 17076 42708 17088
rect 42760 17076 42766 17128
rect 42978 17116 42984 17128
rect 42939 17088 42984 17116
rect 42978 17076 42984 17088
rect 43036 17076 43042 17128
rect 40310 17048 40316 17060
rect 40052 17020 40316 17048
rect 40310 17008 40316 17020
rect 40368 17048 40374 17060
rect 41230 17048 41236 17060
rect 40368 17020 41236 17048
rect 40368 17008 40374 17020
rect 41230 17008 41236 17020
rect 41288 17008 41294 17060
rect 46934 16980 46940 16992
rect 46895 16952 46940 16980
rect 46934 16940 46940 16952
rect 46992 16940 46998 16992
rect 47762 16980 47768 16992
rect 47723 16952 47768 16980
rect 47762 16940 47768 16952
rect 47820 16940 47826 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 2314 16736 2320 16788
rect 2372 16776 2378 16788
rect 2501 16779 2559 16785
rect 2501 16776 2513 16779
rect 2372 16748 2513 16776
rect 2372 16736 2378 16748
rect 2501 16745 2513 16748
rect 2547 16745 2559 16779
rect 39850 16776 39856 16788
rect 39811 16748 39856 16776
rect 2501 16739 2559 16745
rect 39850 16736 39856 16748
rect 39908 16736 39914 16788
rect 40954 16640 40960 16652
rect 40052 16612 40960 16640
rect 2406 16582 2412 16594
rect 2367 16554 2412 16582
rect 2406 16542 2412 16554
rect 2464 16542 2470 16594
rect 40052 16581 40080 16612
rect 40954 16600 40960 16612
rect 41012 16600 41018 16652
rect 46293 16643 46351 16649
rect 46293 16609 46305 16643
rect 46339 16640 46351 16643
rect 47762 16640 47768 16652
rect 46339 16612 47768 16640
rect 46339 16609 46351 16612
rect 46293 16603 46351 16609
rect 47762 16600 47768 16612
rect 47820 16600 47826 16652
rect 48130 16640 48136 16652
rect 48091 16612 48136 16640
rect 48130 16600 48136 16612
rect 48188 16600 48194 16652
rect 40037 16575 40095 16581
rect 40037 16541 40049 16575
rect 40083 16574 40095 16575
rect 40313 16575 40371 16581
rect 40083 16546 40117 16574
rect 40083 16541 40095 16546
rect 40037 16535 40095 16541
rect 40313 16541 40325 16575
rect 40359 16572 40371 16575
rect 40402 16572 40408 16584
rect 40359 16544 40408 16572
rect 40359 16541 40371 16544
rect 40313 16535 40371 16541
rect 40402 16532 40408 16544
rect 40460 16532 40466 16584
rect 46477 16507 46535 16513
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 46934 16504 46940 16516
rect 46523 16476 46940 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 46934 16464 46940 16476
rect 46992 16464 46998 16516
rect 40218 16436 40224 16448
rect 40179 16408 40224 16436
rect 40218 16396 40224 16408
rect 40276 16396 40282 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 2130 15444 2136 15496
rect 2188 15484 2194 15496
rect 2317 15487 2375 15493
rect 2317 15484 2329 15487
rect 2188 15456 2329 15484
rect 2188 15444 2194 15456
rect 2317 15453 2329 15456
rect 2363 15453 2375 15487
rect 47670 15484 47676 15496
rect 47631 15456 47676 15484
rect 2317 15447 2375 15453
rect 47670 15444 47676 15456
rect 47728 15444 47734 15496
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 47578 15008 47584 15020
rect 47539 14980 47584 15008
rect 47578 14968 47584 14980
rect 47636 14968 47642 15020
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14940 2375 14943
rect 2590 14940 2596 14952
rect 2363 14912 2596 14940
rect 2363 14909 2375 14912
rect 2317 14903 2375 14909
rect 2590 14900 2596 14912
rect 2648 14900 2654 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 46474 14764 46480 14816
rect 46532 14804 46538 14816
rect 47673 14807 47731 14813
rect 47673 14804 47685 14807
rect 46532 14776 47685 14804
rect 46532 14764 46538 14776
rect 47673 14773 47685 14776
rect 47719 14773 47731 14807
rect 47673 14767 47731 14773
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 2590 14600 2596 14612
rect 2551 14572 2596 14600
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 47670 14532 47676 14544
rect 46308 14504 47676 14532
rect 8570 14464 8576 14476
rect 1872 14436 8576 14464
rect 1872 14405 1900 14436
rect 8570 14424 8576 14436
rect 8628 14464 8634 14476
rect 9214 14464 9220 14476
rect 8628 14436 9220 14464
rect 8628 14424 8634 14436
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 46308 14473 46336 14504
rect 47670 14492 47676 14504
rect 47728 14492 47734 14544
rect 46293 14467 46351 14473
rect 46293 14433 46305 14467
rect 46339 14433 46351 14467
rect 46474 14464 46480 14476
rect 46435 14436 46480 14464
rect 46293 14427 46351 14433
rect 46474 14424 46480 14436
rect 46532 14424 46538 14476
rect 48130 14464 48136 14476
rect 48091 14436 48136 14464
rect 48130 14424 48136 14436
rect 48188 14424 48194 14476
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14365 1915 14399
rect 2498 14396 2504 14408
rect 2459 14368 2504 14396
rect 1857 14359 1915 14365
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 2130 14288 2136 14340
rect 2188 14328 2194 14340
rect 3988 14328 4016 14359
rect 2188 14300 4016 14328
rect 2188 14288 2194 14300
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 2314 14260 2320 14272
rect 1995 14232 2320 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 2314 13988 2320 14000
rect 2275 13960 2320 13988
rect 2314 13948 2320 13960
rect 2372 13948 2378 14000
rect 2130 13920 2136 13932
rect 2091 13892 2136 13920
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 2774 13852 2780 13864
rect 2735 13824 2780 13852
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 46658 13744 46664 13796
rect 46716 13784 46722 13796
rect 47118 13784 47124 13796
rect 46716 13756 47124 13784
rect 46716 13744 46722 13756
rect 47118 13744 47124 13756
rect 47176 13744 47182 13796
rect 47762 13716 47768 13728
rect 47723 13688 47768 13716
rect 47762 13676 47768 13688
rect 47820 13676 47826 13728
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 46293 13379 46351 13385
rect 46293 13345 46305 13379
rect 46339 13376 46351 13379
rect 47762 13376 47768 13388
rect 46339 13348 47768 13376
rect 46339 13345 46351 13348
rect 46293 13339 46351 13345
rect 47762 13336 47768 13348
rect 47820 13336 47826 13388
rect 48130 13376 48136 13388
rect 48091 13348 48136 13376
rect 48130 13336 48136 13348
rect 48188 13336 48194 13388
rect 46477 13243 46535 13249
rect 46477 13209 46489 13243
rect 46523 13240 46535 13243
rect 47670 13240 47676 13252
rect 46523 13212 47676 13240
rect 46523 13209 46535 13212
rect 46477 13203 46535 13209
rect 47670 13200 47676 13212
rect 47728 13200 47734 13252
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 47670 12968 47676 12980
rect 47631 12940 47676 12968
rect 47670 12928 47676 12940
rect 47728 12928 47734 12980
rect 46201 12835 46259 12841
rect 46201 12801 46213 12835
rect 46247 12832 46259 12835
rect 46658 12832 46664 12844
rect 46247 12804 46664 12832
rect 46247 12801 46259 12804
rect 46201 12795 46259 12801
rect 46658 12792 46664 12804
rect 46716 12792 46722 12844
rect 47578 12832 47584 12844
rect 47539 12804 47584 12832
rect 47578 12792 47584 12804
rect 47636 12792 47642 12844
rect 46293 12631 46351 12637
rect 46293 12597 46305 12631
rect 46339 12628 46351 12631
rect 46474 12628 46480 12640
rect 46339 12600 46480 12628
rect 46339 12597 46351 12600
rect 46293 12591 46351 12597
rect 46474 12588 46480 12600
rect 46532 12588 46538 12640
rect 47026 12628 47032 12640
rect 46987 12600 47032 12628
rect 47026 12588 47032 12600
rect 47084 12588 47090 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 47026 12356 47032 12368
rect 46308 12328 47032 12356
rect 46308 12297 46336 12328
rect 47026 12316 47032 12328
rect 47084 12316 47090 12368
rect 46293 12291 46351 12297
rect 46293 12257 46305 12291
rect 46339 12257 46351 12291
rect 46474 12288 46480 12300
rect 46435 12260 46480 12288
rect 46293 12251 46351 12257
rect 46474 12248 46480 12260
rect 46532 12248 46538 12300
rect 48130 12288 48136 12300
rect 48091 12260 48136 12288
rect 48130 12248 48136 12260
rect 48188 12248 48194 12300
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 2317 12223 2375 12229
rect 2317 12220 2329 12223
rect 2096 12192 2329 12220
rect 2096 12180 2102 12192
rect 2317 12189 2329 12192
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 2038 11744 2044 11756
rect 1999 11716 2044 11744
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 18414 11704 18420 11756
rect 18472 11744 18478 11756
rect 41414 11744 41420 11756
rect 18472 11716 41420 11744
rect 18472 11704 18478 11716
rect 41414 11704 41420 11716
rect 41472 11744 41478 11756
rect 46753 11747 46811 11753
rect 46753 11744 46765 11747
rect 41472 11716 46765 11744
rect 41472 11704 41478 11716
rect 46753 11713 46765 11716
rect 46799 11713 46811 11747
rect 46753 11707 46811 11713
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2774 11676 2780 11688
rect 2735 11648 2780 11676
rect 2774 11636 2780 11648
rect 2832 11636 2838 11688
rect 46474 11500 46480 11552
rect 46532 11540 46538 11552
rect 46845 11543 46903 11549
rect 46845 11540 46857 11543
rect 46532 11512 46857 11540
rect 46532 11500 46538 11512
rect 46845 11509 46857 11512
rect 46891 11509 46903 11543
rect 47762 11540 47768 11552
rect 47723 11512 47768 11540
rect 46845 11503 46903 11509
rect 47762 11500 47768 11512
rect 47820 11500 47826 11552
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 2280 11308 2421 11336
rect 2280 11296 2286 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2409 11299 2467 11305
rect 47762 11268 47768 11280
rect 46308 11240 47768 11268
rect 46308 11209 46336 11240
rect 47762 11228 47768 11240
rect 47820 11228 47826 11280
rect 46293 11203 46351 11209
rect 46293 11169 46305 11203
rect 46339 11169 46351 11203
rect 46474 11200 46480 11212
rect 46435 11172 46480 11200
rect 46293 11163 46351 11169
rect 46474 11160 46480 11172
rect 46532 11160 46538 11212
rect 46842 11200 46848 11212
rect 46803 11172 46848 11200
rect 46842 11160 46848 11172
rect 46900 11160 46906 11212
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2866 11132 2872 11144
rect 2363 11104 2872 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3142 11132 3148 11144
rect 3103 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 3142 10724 3148 10736
rect 2148 10696 3148 10724
rect 2148 10665 2176 10696
rect 3142 10684 3148 10696
rect 3200 10684 3206 10736
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 2314 10588 2320 10600
rect 2275 10560 2320 10588
rect 2314 10548 2320 10560
rect 2372 10548 2378 10600
rect 3694 10588 3700 10600
rect 3655 10560 3700 10588
rect 3694 10548 3700 10560
rect 3752 10548 3758 10600
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 22094 10452 22100 10464
rect 5500 10424 22100 10452
rect 5500 10412 5506 10424
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 2225 10251 2283 10257
rect 2225 10217 2237 10251
rect 2271 10248 2283 10251
rect 2314 10248 2320 10260
rect 2271 10220 2320 10248
rect 2271 10217 2283 10220
rect 2225 10211 2283 10217
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 2832 10016 2973 10044
rect 2832 10004 2838 10016
rect 2961 10013 2973 10016
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10044 3847 10047
rect 5442 10044 5448 10056
rect 3835 10016 5448 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10044 19763 10047
rect 19978 10044 19984 10056
rect 19751 10016 19984 10044
rect 19751 10013 19763 10016
rect 19705 10007 19763 10013
rect 19978 10004 19984 10016
rect 20036 10044 20042 10056
rect 26421 10047 26479 10053
rect 26421 10044 26433 10047
rect 20036 10016 26433 10044
rect 20036 10004 20042 10016
rect 26421 10013 26433 10016
rect 26467 10013 26479 10047
rect 26421 10007 26479 10013
rect 20070 9976 20076 9988
rect 20031 9948 20076 9976
rect 20070 9936 20076 9948
rect 20128 9936 20134 9988
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3016 9880 3893 9908
rect 3016 9868 3022 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 26513 9911 26571 9917
rect 26513 9877 26525 9911
rect 26559 9908 26571 9911
rect 27154 9908 27160 9920
rect 26559 9880 27160 9908
rect 26559 9877 26571 9880
rect 26513 9871 26571 9877
rect 27154 9868 27160 9880
rect 27212 9868 27218 9920
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 2958 9636 2964 9648
rect 2919 9608 2964 9636
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 2130 9568 2136 9580
rect 2043 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2774 9568 2780 9580
rect 2735 9540 2780 9568
rect 2774 9528 2780 9540
rect 2832 9528 2838 9580
rect 2148 9432 2176 9528
rect 3234 9500 3240 9512
rect 3195 9472 3240 9500
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 7190 9432 7196 9444
rect 2148 9404 7196 9432
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 2314 9364 2320 9376
rect 2271 9336 2320 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 2188 8928 2329 8956
rect 2188 8916 2194 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 45830 8576 45836 8628
rect 45888 8616 45894 8628
rect 48041 8619 48099 8625
rect 48041 8616 48053 8619
rect 45888 8588 48053 8616
rect 45888 8576 45894 8588
rect 48041 8585 48053 8588
rect 48087 8585 48099 8619
rect 48041 8579 48099 8585
rect 2314 8548 2320 8560
rect 2275 8520 2320 8548
rect 2314 8508 2320 8520
rect 2372 8508 2378 8560
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 47946 8480 47952 8492
rect 47907 8452 47952 8480
rect 47946 8440 47952 8452
rect 48004 8440 48010 8492
rect 2866 8412 2872 8424
rect 2827 8384 2872 8412
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 2222 7896 2228 7948
rect 2280 7936 2286 7948
rect 2280 7908 2820 7936
rect 2280 7896 2286 7908
rect 2130 7828 2136 7880
rect 2188 7868 2194 7880
rect 2792 7877 2820 7908
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 2188 7840 2329 7868
rect 2188 7828 2194 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2958 7868 2964 7880
rect 2823 7840 2964 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2869 7735 2927 7741
rect 2869 7732 2881 7735
rect 2372 7704 2881 7732
rect 2372 7692 2378 7704
rect 2869 7701 2881 7704
rect 2915 7701 2927 7735
rect 2869 7695 2927 7701
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 2314 7460 2320 7472
rect 2275 7432 2320 7460
rect 2314 7420 2320 7432
rect 2372 7420 2378 7472
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 47578 7392 47584 7404
rect 47539 7364 47584 7392
rect 47578 7352 47584 7364
rect 47636 7352 47642 7404
rect 2774 7324 2780 7336
rect 2735 7296 2780 7324
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 1670 7188 1676 7200
rect 1631 7160 1676 7188
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 47670 7188 47676 7200
rect 47631 7160 47676 7188
rect 47670 7148 47676 7160
rect 47728 7148 47734 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 46477 6851 46535 6857
rect 46477 6817 46489 6851
rect 46523 6848 46535 6851
rect 47670 6848 47676 6860
rect 46523 6820 47676 6848
rect 46523 6817 46535 6820
rect 46477 6811 46535 6817
rect 47670 6808 47676 6820
rect 47728 6808 47734 6860
rect 48130 6848 48136 6860
rect 48091 6820 48136 6848
rect 48130 6808 48136 6820
rect 48188 6808 48194 6860
rect 2406 6780 2412 6792
rect 2367 6752 2412 6780
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 46293 6783 46351 6789
rect 46293 6749 46305 6783
rect 46339 6749 46351 6783
rect 46293 6743 46351 6749
rect 46308 6712 46336 6743
rect 47762 6712 47768 6724
rect 46308 6684 47768 6712
rect 47762 6672 47768 6684
rect 47820 6672 47826 6724
rect 2314 6604 2320 6656
rect 2372 6644 2378 6656
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 2372 6616 2513 6644
rect 2372 6604 2378 6616
rect 2501 6613 2513 6616
rect 2547 6613 2559 6647
rect 2501 6607 2559 6613
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 2314 6372 2320 6384
rect 2275 6344 2320 6372
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 47486 6372 47492 6384
rect 46216 6344 47492 6372
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1728 6276 2145 6304
rect 1728 6264 1734 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 45554 6264 45560 6316
rect 45612 6304 45618 6316
rect 46216 6313 46244 6344
rect 47486 6332 47492 6344
rect 47544 6332 47550 6384
rect 46201 6307 46259 6313
rect 46201 6304 46213 6307
rect 45612 6276 46213 6304
rect 45612 6264 45618 6276
rect 46201 6273 46213 6276
rect 46247 6273 46259 6307
rect 46201 6267 46259 6273
rect 46658 6264 46664 6316
rect 46716 6304 46722 6316
rect 46845 6307 46903 6313
rect 46845 6304 46857 6307
rect 46716 6276 46857 6304
rect 46716 6264 46722 6276
rect 46845 6273 46857 6276
rect 46891 6273 46903 6307
rect 47762 6304 47768 6316
rect 47723 6276 47768 6304
rect 46845 6267 46903 6273
rect 47762 6264 47768 6276
rect 47820 6264 47826 6316
rect 2774 6236 2780 6248
rect 2735 6208 2780 6236
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 46290 6100 46296 6112
rect 46251 6072 46296 6100
rect 46290 6060 46296 6072
rect 46348 6060 46354 6112
rect 46934 6100 46940 6112
rect 46895 6072 46940 6100
rect 46934 6060 46940 6072
rect 46992 6060 46998 6112
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 1949 5695 2007 5701
rect 1949 5692 1961 5695
rect 1728 5664 1961 5692
rect 1728 5652 1734 5664
rect 1949 5661 1961 5664
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2406 5652 2412 5704
rect 2464 5692 2470 5704
rect 2593 5695 2651 5701
rect 2593 5692 2605 5695
rect 2464 5664 2605 5692
rect 2464 5652 2470 5664
rect 2593 5661 2605 5664
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 17218 5692 17224 5704
rect 3835 5664 17224 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 17218 5652 17224 5664
rect 17276 5692 17282 5704
rect 17862 5692 17868 5704
rect 17276 5664 17868 5692
rect 17276 5652 17282 5664
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 45646 5692 45652 5704
rect 45607 5664 45652 5692
rect 45646 5652 45652 5664
rect 45704 5652 45710 5704
rect 45830 5652 45836 5704
rect 45888 5692 45894 5704
rect 46293 5695 46351 5701
rect 46293 5692 46305 5695
rect 45888 5664 46305 5692
rect 45888 5652 45894 5664
rect 46293 5661 46305 5664
rect 46339 5661 46351 5695
rect 46293 5655 46351 5661
rect 45741 5627 45799 5633
rect 45741 5593 45753 5627
rect 45787 5624 45799 5627
rect 46477 5627 46535 5633
rect 46477 5624 46489 5627
rect 45787 5596 46489 5624
rect 45787 5593 45799 5596
rect 45741 5587 45799 5593
rect 46477 5593 46489 5596
rect 46523 5593 46535 5627
rect 46477 5587 46535 5593
rect 48133 5627 48191 5633
rect 48133 5593 48145 5627
rect 48179 5624 48191 5627
rect 48222 5624 48228 5636
rect 48179 5596 48228 5624
rect 48179 5593 48191 5596
rect 48133 5587 48191 5593
rect 48222 5584 48228 5596
rect 48280 5584 48286 5636
rect 3878 5556 3884 5568
rect 3839 5528 3884 5556
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 4062 5352 4068 5364
rect 2832 5324 4068 5352
rect 2832 5312 2838 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 2593 5287 2651 5293
rect 2593 5253 2605 5287
rect 2639 5284 2651 5287
rect 3878 5284 3884 5296
rect 2639 5256 3884 5284
rect 2639 5253 2651 5256
rect 2593 5247 2651 5253
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 45373 5287 45431 5293
rect 45373 5253 45385 5287
rect 45419 5284 45431 5287
rect 46290 5284 46296 5296
rect 45419 5256 46296 5284
rect 45419 5253 45431 5256
rect 45373 5247 45431 5253
rect 46290 5244 46296 5256
rect 46348 5244 46354 5296
rect 2406 5216 2412 5228
rect 2367 5188 2412 5216
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2866 5148 2872 5160
rect 2827 5120 2872 5148
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 44729 5151 44787 5157
rect 44729 5117 44741 5151
rect 44775 5148 44787 5151
rect 45189 5151 45247 5157
rect 45189 5148 45201 5151
rect 44775 5120 45201 5148
rect 44775 5117 44787 5120
rect 44729 5111 44787 5117
rect 45189 5117 45201 5120
rect 45235 5117 45247 5151
rect 46842 5148 46848 5160
rect 46803 5120 46848 5148
rect 45189 5111 45247 5117
rect 46842 5108 46848 5120
rect 46900 5108 46906 5160
rect 1946 5012 1952 5024
rect 1907 4984 1952 5012
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 46290 4972 46296 5024
rect 46348 5012 46354 5024
rect 47765 5015 47823 5021
rect 47765 5012 47777 5015
rect 46348 4984 47777 5012
rect 46348 4972 46354 4984
rect 47765 4981 47777 4984
rect 47811 4981 47823 5015
rect 47765 4975 47823 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 8018 4808 8024 4820
rect 2976 4780 8024 4808
rect 2866 4672 2872 4684
rect 1688 4644 2872 4672
rect 1688 4613 1716 4644
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2774 4604 2780 4616
rect 2363 4576 2780 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 2976 4613 3004 4780
rect 8018 4768 8024 4780
rect 8076 4808 8082 4820
rect 14090 4808 14096 4820
rect 8076 4780 14096 4808
rect 8076 4768 8082 4780
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 44453 4811 44511 4817
rect 44453 4777 44465 4811
rect 44499 4808 44511 4811
rect 45830 4808 45836 4820
rect 44499 4780 45836 4808
rect 44499 4777 44511 4780
rect 44453 4771 44511 4777
rect 45830 4768 45836 4780
rect 45888 4768 45894 4820
rect 46290 4672 46296 4684
rect 46251 4644 46296 4672
rect 46290 4632 46296 4644
rect 46348 4632 46354 4684
rect 46477 4675 46535 4681
rect 46477 4641 46489 4675
rect 46523 4672 46535 4675
rect 46934 4672 46940 4684
rect 46523 4644 46940 4672
rect 46523 4641 46535 4644
rect 46477 4635 46535 4641
rect 46934 4632 46940 4644
rect 46992 4632 46998 4684
rect 48130 4672 48136 4684
rect 48091 4644 48136 4672
rect 48130 4632 48136 4644
rect 48188 4632 48194 4684
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4706 4604 4712 4616
rect 4479 4576 4712 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4536 1823 4539
rect 3970 4536 3976 4548
rect 1811 4508 3976 4536
rect 1811 4505 1823 4508
rect 1765 4499 1823 4505
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 4522 4496 4528 4548
rect 4580 4536 4586 4548
rect 4908 4536 4936 4567
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 6144 4576 6377 4604
rect 6144 4564 6150 4576
rect 6365 4573 6377 4576
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7800 4576 8033 4604
rect 7800 4564 7806 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 9030 4604 9036 4616
rect 8987 4576 9036 4604
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 17310 4564 17316 4616
rect 17368 4604 17374 4616
rect 19245 4607 19303 4613
rect 19245 4604 19257 4607
rect 17368 4576 19257 4604
rect 17368 4564 17374 4576
rect 19245 4573 19257 4576
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4604 19947 4607
rect 20070 4604 20076 4616
rect 19935 4576 20076 4604
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 42334 4604 42340 4616
rect 42295 4576 42340 4604
rect 42334 4564 42340 4576
rect 42392 4564 42398 4616
rect 45281 4607 45339 4613
rect 45281 4573 45293 4607
rect 45327 4604 45339 4607
rect 46198 4604 46204 4616
rect 45327 4576 46204 4604
rect 45327 4573 45339 4576
rect 45281 4567 45339 4573
rect 46198 4564 46204 4576
rect 46256 4564 46262 4616
rect 20438 4536 20444 4548
rect 4580 4508 20444 4536
rect 4580 4496 4586 4508
rect 20438 4496 20444 4508
rect 20496 4496 20502 4548
rect 2406 4468 2412 4480
rect 2367 4440 2412 4468
rect 2406 4428 2412 4440
rect 2464 4428 2470 4480
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 4982 4468 4988 4480
rect 4943 4440 4988 4468
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 8570 4428 8576 4480
rect 8628 4468 8634 4480
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 8628 4440 9045 4468
rect 8628 4428 8634 4440
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 19334 4468 19340 4480
rect 19295 4440 19340 4468
rect 9033 4431 9091 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 19978 4468 19984 4480
rect 19939 4440 19984 4468
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 45370 4468 45376 4480
rect 45331 4440 45376 4468
rect 45370 4428 45376 4440
rect 45428 4428 45434 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 41506 4264 41512 4276
rect 39868 4236 41512 4264
rect 1486 4128 1492 4140
rect 1447 4100 1492 4128
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2133 4131 2191 4137
rect 2133 4128 2145 4131
rect 2004 4100 2145 4128
rect 2004 4088 2010 4100
rect 2133 4097 2145 4100
rect 2179 4097 2191 4131
rect 4522 4128 4528 4140
rect 4483 4100 4528 4128
rect 2133 4091 2191 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 6362 4128 6368 4140
rect 6323 4100 6368 4128
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7190 4128 7196 4140
rect 7147 4100 7196 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7742 4128 7748 4140
rect 7703 4100 7748 4128
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 22094 4128 22100 4140
rect 22055 4100 22100 4128
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 25409 4131 25467 4137
rect 25409 4097 25421 4131
rect 25455 4097 25467 4131
rect 38654 4128 38660 4140
rect 38567 4100 38660 4128
rect 25409 4091 25467 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 3050 4060 3056 4072
rect 2363 4032 3056 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 7929 4063 7987 4069
rect 3200 4032 3245 4060
rect 3200 4020 3206 4032
rect 7929 4029 7941 4063
rect 7975 4060 7987 4063
rect 8570 4060 8576 4072
rect 7975 4032 8576 4060
rect 7975 4029 7987 4032
rect 7929 4023 7987 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 8665 4063 8723 4069
rect 8665 4029 8677 4063
rect 8711 4029 8723 4063
rect 12342 4060 12348 4072
rect 12303 4032 12348 4060
rect 8665 4023 8723 4029
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 8680 3992 8708 4023
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 12802 4060 12808 4072
rect 12575 4032 12808 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12894 4020 12900 4072
rect 12952 4060 12958 4072
rect 18233 4063 18291 4069
rect 12952 4032 12997 4060
rect 12952 4020 12958 4032
rect 18233 4029 18245 4063
rect 18279 4060 18291 4063
rect 18693 4063 18751 4069
rect 18693 4060 18705 4063
rect 18279 4032 18705 4060
rect 18279 4029 18291 4032
rect 18233 4023 18291 4029
rect 18693 4029 18705 4032
rect 18739 4029 18751 4063
rect 18693 4023 18751 4029
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4060 18935 4063
rect 19334 4060 19340 4072
rect 18923 4032 19340 4060
rect 18923 4029 18935 4032
rect 18877 4023 18935 4029
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19484 4032 19529 4060
rect 19484 4020 19490 4032
rect 7156 3964 8708 3992
rect 7156 3952 7162 3964
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 25424 3992 25452 4091
rect 38654 4088 38660 4100
rect 38712 4128 38718 4140
rect 39868 4128 39896 4236
rect 41506 4224 41512 4236
rect 41564 4224 41570 4276
rect 45554 4264 45560 4276
rect 45204 4236 45560 4264
rect 38712 4100 39896 4128
rect 39960 4168 40172 4196
rect 38712 4088 38718 4100
rect 39960 4060 39988 4168
rect 40037 4131 40095 4137
rect 40037 4097 40049 4131
rect 40083 4097 40095 4131
rect 40037 4091 40095 4097
rect 26206 4032 39988 4060
rect 26206 3992 26234 4032
rect 9272 3964 26234 3992
rect 9272 3952 9278 3964
rect 38562 3952 38568 4004
rect 38620 3992 38626 4004
rect 39485 3995 39543 4001
rect 39485 3992 39497 3995
rect 38620 3964 39497 3992
rect 38620 3952 38626 3964
rect 39485 3961 39497 3964
rect 39531 3961 39543 3995
rect 40052 3992 40080 4091
rect 40144 4060 40172 4168
rect 41966 4156 41972 4208
rect 42024 4196 42030 4208
rect 42024 4168 42656 4196
rect 42024 4156 42030 4168
rect 40770 4128 40776 4140
rect 40731 4100 40776 4128
rect 40770 4088 40776 4100
rect 40828 4088 40834 4140
rect 41386 4106 41644 4134
rect 41386 4060 41414 4106
rect 40144 4032 41414 4060
rect 41616 4060 41644 4106
rect 41693 4131 41751 4137
rect 41693 4097 41705 4131
rect 41739 4128 41751 4131
rect 42518 4128 42524 4140
rect 41739 4100 42524 4128
rect 41739 4097 41751 4100
rect 41693 4091 41751 4097
rect 42518 4088 42524 4100
rect 42576 4088 42582 4140
rect 42628 4128 42656 4168
rect 43456 4168 43668 4196
rect 43456 4128 43484 4168
rect 42628 4100 43484 4128
rect 43533 4131 43591 4137
rect 43533 4097 43545 4131
rect 43579 4097 43591 4131
rect 43640 4128 43668 4168
rect 45204 4128 45232 4236
rect 45554 4224 45560 4236
rect 45612 4224 45618 4276
rect 45370 4196 45376 4208
rect 45331 4168 45376 4196
rect 45370 4156 45376 4168
rect 45428 4156 45434 4208
rect 43640 4100 45232 4128
rect 43533 4091 43591 4097
rect 43548 4060 43576 4091
rect 41616 4032 43576 4060
rect 45189 4063 45247 4069
rect 45189 4029 45201 4063
rect 45235 4029 45247 4063
rect 47026 4060 47032 4072
rect 46987 4032 47032 4060
rect 45189 4023 45247 4029
rect 41414 3992 41420 4004
rect 40052 3964 41420 3992
rect 39485 3955 39543 3961
rect 41414 3952 41420 3964
rect 41472 3952 41478 4004
rect 41506 3952 41512 4004
rect 41564 3992 41570 4004
rect 45204 3992 45232 4023
rect 47026 4020 47032 4032
rect 47084 4020 47090 4072
rect 47765 3995 47823 4001
rect 47765 3992 47777 3995
rect 41564 3964 44864 3992
rect 45204 3964 47777 3992
rect 41564 3952 41570 3964
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5810 3924 5816 3936
rect 5771 3896 5816 3924
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 6328 3896 6469 3924
rect 6328 3884 6334 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 6457 3887 6515 3893
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 9122 3924 9128 3936
rect 7239 3896 9128 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 10689 3927 10747 3933
rect 10689 3924 10701 3927
rect 10468 3896 10701 3924
rect 10468 3884 10474 3896
rect 10689 3893 10701 3896
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17184 3896 17417 3924
rect 17184 3884 17190 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 22186 3924 22192 3936
rect 22147 3896 22192 3924
rect 17405 3887 17463 3893
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 25498 3924 25504 3936
rect 25459 3896 25504 3924
rect 25498 3884 25504 3896
rect 25556 3884 25562 3936
rect 38746 3924 38752 3936
rect 38707 3896 38752 3924
rect 38746 3884 38752 3896
rect 38804 3884 38810 3936
rect 40034 3884 40040 3936
rect 40092 3924 40098 3936
rect 40129 3927 40187 3933
rect 40129 3924 40141 3927
rect 40092 3896 40141 3924
rect 40092 3884 40098 3896
rect 40129 3893 40141 3896
rect 40175 3893 40187 3927
rect 40862 3924 40868 3936
rect 40823 3896 40868 3924
rect 40129 3887 40187 3893
rect 40862 3884 40868 3896
rect 40920 3884 40926 3936
rect 41782 3924 41788 3936
rect 41743 3896 41788 3924
rect 41782 3884 41788 3896
rect 41840 3884 41846 3936
rect 42150 3884 42156 3936
rect 42208 3924 42214 3936
rect 42613 3927 42671 3933
rect 42613 3924 42625 3927
rect 42208 3896 42625 3924
rect 42208 3884 42214 3896
rect 42613 3893 42625 3896
rect 42659 3893 42671 3927
rect 43622 3924 43628 3936
rect 43583 3896 43628 3924
rect 42613 3887 42671 3893
rect 43622 3884 43628 3896
rect 43680 3884 43686 3936
rect 44361 3927 44419 3933
rect 44361 3893 44373 3927
rect 44407 3924 44419 3927
rect 44726 3924 44732 3936
rect 44407 3896 44732 3924
rect 44407 3893 44419 3896
rect 44361 3887 44419 3893
rect 44726 3884 44732 3896
rect 44784 3884 44790 3936
rect 44836 3924 44864 3964
rect 47765 3961 47777 3964
rect 47811 3961 47823 3995
rect 47765 3955 47823 3961
rect 47578 3924 47584 3936
rect 44836 3896 47584 3924
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 12802 3720 12808 3732
rect 12763 3692 12808 3720
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14148 3692 25728 3720
rect 14148 3680 14154 3692
rect 1486 3612 1492 3664
rect 1544 3652 1550 3664
rect 1544 3624 6914 3652
rect 1544 3612 1550 3624
rect 1578 3584 1584 3596
rect 1539 3556 1584 3584
rect 1578 3544 1584 3556
rect 1636 3544 1642 3596
rect 1854 3584 1860 3596
rect 1815 3556 1860 3584
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 3970 3584 3976 3596
rect 3931 3556 3976 3584
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4120 3556 4261 3584
rect 4120 3544 4126 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 4249 3547 4307 3553
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6270 3584 6276 3596
rect 6231 3556 6276 3584
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 6549 3587 6607 3593
rect 6549 3584 6561 3587
rect 6512 3556 6561 3584
rect 6512 3544 6518 3556
rect 6549 3553 6561 3556
rect 6595 3553 6607 3587
rect 6886 3584 6914 3624
rect 7190 3612 7196 3664
rect 7248 3652 7254 3664
rect 7248 3624 16574 3652
rect 7248 3612 7254 3624
rect 9398 3584 9404 3596
rect 6886 3556 9404 3584
rect 6549 3547 6607 3553
rect 9398 3544 9404 3556
rect 9456 3584 9462 3596
rect 10410 3584 10416 3596
rect 9456 3556 9904 3584
rect 10371 3556 10416 3584
rect 9456 3544 9462 3556
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 3786 3516 3792 3528
rect 3747 3488 3792 3516
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3516 8999 3519
rect 9674 3516 9680 3528
rect 8987 3488 9680 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 7834 3408 7840 3460
rect 7892 3448 7898 3460
rect 9784 3448 9812 3479
rect 7892 3420 9812 3448
rect 7892 3408 7898 3420
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8076 3352 9045 3380
rect 8076 3340 8082 3352
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9876 3380 9904 3556
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 16546 3584 16574 3624
rect 17862 3612 17868 3664
rect 17920 3652 17926 3664
rect 25590 3652 25596 3664
rect 17920 3624 25596 3652
rect 17920 3612 17926 3624
rect 25590 3612 25596 3624
rect 25648 3612 25654 3664
rect 20070 3584 20076 3596
rect 16546 3556 20076 3584
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 10597 3451 10655 3457
rect 10597 3417 10609 3451
rect 10643 3448 10655 3451
rect 10686 3448 10692 3460
rect 10643 3420 10692 3448
rect 10643 3417 10655 3420
rect 10597 3411 10655 3417
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 12728 3380 12756 3479
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13504 3488 13553 3516
rect 13504 3476 13510 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 13541 3479 13599 3485
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 17880 3525 17908 3556
rect 20070 3544 20076 3556
rect 20128 3544 20134 3596
rect 25498 3584 25504 3596
rect 25459 3556 25504 3584
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 25700 3584 25728 3692
rect 25774 3680 25780 3732
rect 25832 3720 25838 3732
rect 25832 3692 28304 3720
rect 25832 3680 25838 3692
rect 28166 3652 28172 3664
rect 26206 3624 28172 3652
rect 26206 3584 26234 3624
rect 28166 3612 28172 3624
rect 28224 3612 28230 3664
rect 25700 3556 26234 3584
rect 26697 3587 26755 3593
rect 26697 3553 26709 3587
rect 26743 3553 26755 3587
rect 26697 3547 26755 3553
rect 28276 3584 28304 3692
rect 41874 3680 41880 3732
rect 41932 3720 41938 3732
rect 45646 3720 45652 3732
rect 41932 3692 42656 3720
rect 41932 3680 41938 3692
rect 28350 3612 28356 3664
rect 28408 3652 28414 3664
rect 28408 3624 40724 3652
rect 28408 3612 28414 3624
rect 40034 3584 40040 3596
rect 28276 3556 32260 3584
rect 39995 3556 40040 3584
rect 17221 3519 17279 3525
rect 17221 3485 17233 3519
rect 17267 3516 17279 3519
rect 17865 3519 17923 3525
rect 17267 3488 17816 3516
rect 17267 3485 17279 3488
rect 17221 3479 17279 3485
rect 9876 3352 12756 3380
rect 9033 3343 9091 3349
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13688 3352 14197 3380
rect 13688 3340 13694 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 14185 3343 14243 3349
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 17788 3380 17816 3488
rect 17865 3485 17877 3519
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 18739 3488 19533 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 22002 3476 22008 3528
rect 22060 3516 22066 3528
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 22060 3488 22201 3516
rect 22060 3476 22066 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 25314 3516 25320 3528
rect 25275 3488 25320 3516
rect 22189 3479 22247 3485
rect 25314 3476 25320 3488
rect 25372 3476 25378 3528
rect 17957 3451 18015 3457
rect 17957 3417 17969 3451
rect 18003 3448 18015 3451
rect 19705 3451 19763 3457
rect 19705 3448 19717 3451
rect 18003 3420 19717 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 19705 3417 19717 3420
rect 19751 3417 19763 3451
rect 21358 3448 21364 3460
rect 21319 3420 21364 3448
rect 19705 3411 19763 3417
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 25774 3408 25780 3460
rect 25832 3448 25838 3460
rect 26712 3448 26740 3547
rect 27798 3516 27804 3528
rect 27759 3488 27804 3516
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 28276 3525 28304 3556
rect 28261 3519 28319 3525
rect 28261 3485 28273 3519
rect 28307 3485 28319 3519
rect 28261 3479 28319 3485
rect 31757 3519 31815 3525
rect 31757 3485 31769 3519
rect 31803 3516 31815 3519
rect 32122 3516 32128 3528
rect 31803 3488 32128 3516
rect 31803 3485 31815 3488
rect 31757 3479 31815 3485
rect 32122 3476 32128 3488
rect 32180 3476 32186 3528
rect 32232 3525 32260 3556
rect 40034 3544 40040 3556
rect 40092 3544 40098 3596
rect 40586 3584 40592 3596
rect 40547 3556 40592 3584
rect 40586 3544 40592 3556
rect 40644 3544 40650 3596
rect 40696 3584 40724 3624
rect 41782 3612 41788 3664
rect 41840 3652 41846 3664
rect 41840 3624 42380 3652
rect 41840 3612 41846 3624
rect 41966 3584 41972 3596
rect 40696 3556 41972 3584
rect 41966 3544 41972 3556
rect 42024 3544 42030 3596
rect 42150 3584 42156 3596
rect 42111 3556 42156 3584
rect 42150 3544 42156 3556
rect 42208 3544 42214 3596
rect 42352 3593 42380 3624
rect 42628 3593 42656 3692
rect 43548 3692 45652 3720
rect 42337 3587 42395 3593
rect 42337 3553 42349 3587
rect 42383 3553 42395 3587
rect 42337 3547 42395 3553
rect 42613 3587 42671 3593
rect 42613 3553 42625 3587
rect 42659 3553 42671 3587
rect 42613 3547 42671 3553
rect 32217 3519 32275 3525
rect 32217 3485 32229 3519
rect 32263 3485 32275 3519
rect 32217 3479 32275 3485
rect 39301 3519 39359 3525
rect 39301 3485 39313 3519
rect 39347 3516 39359 3519
rect 39853 3519 39911 3525
rect 39853 3516 39865 3519
rect 39347 3488 39865 3516
rect 39347 3485 39359 3488
rect 39301 3479 39359 3485
rect 39853 3485 39865 3488
rect 39899 3485 39911 3519
rect 39853 3479 39911 3485
rect 25832 3420 26740 3448
rect 28184 3420 35894 3448
rect 25832 3408 25838 3420
rect 18598 3380 18604 3392
rect 17788 3352 18604 3380
rect 18598 3340 18604 3352
rect 18656 3380 18662 3392
rect 28184 3380 28212 3420
rect 28350 3380 28356 3392
rect 18656 3352 28212 3380
rect 28311 3352 28356 3380
rect 18656 3340 18662 3352
rect 28350 3340 28356 3352
rect 28408 3340 28414 3392
rect 32306 3380 32312 3392
rect 32267 3352 32312 3380
rect 32306 3340 32312 3352
rect 32364 3340 32370 3392
rect 35866 3380 35894 3420
rect 38470 3408 38476 3460
rect 38528 3448 38534 3460
rect 43346 3448 43352 3460
rect 38528 3420 43352 3448
rect 38528 3408 38534 3420
rect 43346 3408 43352 3420
rect 43404 3408 43410 3460
rect 43548 3380 43576 3692
rect 45646 3680 45652 3692
rect 45704 3680 45710 3732
rect 46382 3652 46388 3664
rect 45020 3624 46388 3652
rect 45020 3525 45048 3624
rect 46382 3612 46388 3624
rect 46440 3612 46446 3664
rect 46293 3587 46351 3593
rect 46293 3553 46305 3587
rect 46339 3584 46351 3587
rect 47486 3584 47492 3596
rect 46339 3556 47492 3584
rect 46339 3553 46351 3556
rect 46293 3547 46351 3553
rect 47486 3544 47492 3556
rect 47544 3544 47550 3596
rect 47762 3584 47768 3596
rect 47723 3556 47768 3584
rect 47762 3544 47768 3556
rect 47820 3544 47826 3596
rect 45005 3519 45063 3525
rect 45005 3485 45017 3519
rect 45051 3485 45063 3519
rect 45830 3516 45836 3528
rect 45791 3488 45836 3516
rect 45005 3479 45063 3485
rect 45830 3476 45836 3488
rect 45888 3476 45894 3528
rect 46477 3451 46535 3457
rect 46477 3417 46489 3451
rect 46523 3448 46535 3451
rect 47670 3448 47676 3460
rect 46523 3420 47676 3448
rect 46523 3417 46535 3420
rect 46477 3411 46535 3417
rect 47670 3408 47676 3420
rect 47728 3408 47734 3460
rect 35866 3352 43576 3380
rect 45097 3383 45155 3389
rect 45097 3349 45109 3383
rect 45143 3380 45155 3383
rect 45186 3380 45192 3392
rect 45143 3352 45192 3380
rect 45143 3349 45155 3352
rect 45097 3343 45155 3349
rect 45186 3340 45192 3352
rect 45244 3340 45250 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 10686 3176 10692 3188
rect 6886 3148 9260 3176
rect 10647 3148 10692 3176
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 2406 3108 2412 3120
rect 1903 3080 2412 3108
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 4157 3111 4215 3117
rect 4157 3077 4169 3111
rect 4203 3108 4215 3111
rect 4614 3108 4620 3120
rect 4203 3080 4620 3108
rect 4203 3077 4215 3080
rect 4157 3071 4215 3077
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6886 3040 6914 3148
rect 8018 3108 8024 3120
rect 7979 3080 8024 3108
rect 8018 3068 8024 3080
rect 8076 3068 8082 3120
rect 7834 3040 7840 3052
rect 6595 3012 6914 3040
rect 7795 3012 7840 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 9232 3040 9260 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 18874 3176 18880 3188
rect 12728 3148 18880 3176
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 12728 3108 12756 3148
rect 18874 3136 18880 3148
rect 18932 3176 18938 3188
rect 18932 3148 20576 3176
rect 18932 3136 18938 3148
rect 13630 3108 13636 3120
rect 9732 3080 12756 3108
rect 13591 3080 13636 3108
rect 9732 3068 9738 3080
rect 13630 3068 13636 3080
rect 13688 3068 13694 3120
rect 17310 3108 17316 3120
rect 17271 3080 17316 3108
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 19978 3108 19984 3120
rect 19659 3080 19984 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 20548 3108 20576 3148
rect 21358 3136 21364 3188
rect 21416 3176 21422 3188
rect 38470 3176 38476 3188
rect 21416 3148 38476 3176
rect 21416 3136 21422 3148
rect 38470 3136 38476 3148
rect 38528 3136 38534 3188
rect 47670 3176 47676 3188
rect 38580 3148 44496 3176
rect 47631 3148 47676 3176
rect 38580 3108 38608 3148
rect 38746 3108 38752 3120
rect 20548 3080 38608 3108
rect 38707 3080 38752 3108
rect 38746 3068 38752 3080
rect 38804 3068 38810 3120
rect 40862 3068 40868 3120
rect 40920 3108 40926 3120
rect 42613 3111 42671 3117
rect 42613 3108 42625 3111
rect 40920 3080 42625 3108
rect 40920 3068 40926 3080
rect 42613 3077 42625 3080
rect 42659 3077 42671 3111
rect 44468 3108 44496 3148
rect 47670 3136 47676 3148
rect 47728 3136 47734 3188
rect 44468 3080 47624 3108
rect 42613 3071 42671 3077
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 9232 3012 10609 3040
rect 10597 3009 10609 3012
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 2774 2972 2780 2984
rect 2735 2944 2780 2972
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 4706 2972 4712 2984
rect 4019 2944 4712 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 4801 2975 4859 2981
rect 4801 2941 4813 2975
rect 4847 2941 4859 2975
rect 4801 2935 4859 2941
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2941 8539 2975
rect 10612 2972 10640 3003
rect 12342 3000 12348 3052
rect 12400 3040 12406 3052
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 12400 3012 12633 3040
rect 12400 3000 12406 3012
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 13446 3040 13452 3052
rect 13407 3012 13452 3040
rect 12621 3003 12679 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 25314 3000 25320 3052
rect 25372 3040 25378 3052
rect 25593 3043 25651 3049
rect 25593 3040 25605 3043
rect 25372 3012 25605 3040
rect 25372 3000 25378 3012
rect 25593 3009 25605 3012
rect 25639 3009 25651 3043
rect 32122 3040 32128 3052
rect 32083 3012 32128 3040
rect 25593 3003 25651 3009
rect 32122 3000 32128 3012
rect 32180 3000 32186 3052
rect 38562 3040 38568 3052
rect 38523 3012 38568 3040
rect 38562 3000 38568 3012
rect 38620 3000 38626 3052
rect 40770 3040 40776 3052
rect 39960 3012 40776 3040
rect 13078 2972 13084 2984
rect 10612 2944 13084 2972
rect 8481 2935 8539 2941
rect 658 2864 664 2916
rect 716 2904 722 2916
rect 4816 2904 4844 2935
rect 716 2876 4844 2904
rect 716 2864 722 2876
rect 5166 2864 5172 2916
rect 5224 2904 5230 2916
rect 8496 2904 8524 2935
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 13556 2944 13921 2972
rect 13556 2916 13584 2944
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 17589 2975 17647 2981
rect 17589 2972 17601 2975
rect 17460 2944 17601 2972
rect 17460 2932 17466 2944
rect 17589 2941 17601 2944
rect 17635 2941 17647 2975
rect 19426 2972 19432 2984
rect 19387 2944 19432 2972
rect 17589 2935 17647 2941
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 20622 2972 20628 2984
rect 20583 2944 20628 2972
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 22186 2972 22192 2984
rect 22147 2944 22192 2972
rect 22186 2932 22192 2944
rect 22244 2932 22250 2984
rect 22554 2972 22560 2984
rect 22515 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 26421 2975 26479 2981
rect 26421 2941 26433 2975
rect 26467 2972 26479 2975
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26467 2944 26985 2972
rect 26467 2941 26479 2944
rect 26421 2935 26479 2941
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 27154 2972 27160 2984
rect 27115 2944 27160 2972
rect 26973 2935 27031 2941
rect 27154 2932 27160 2944
rect 27212 2932 27218 2984
rect 27246 2932 27252 2984
rect 27304 2972 27310 2984
rect 27433 2975 27491 2981
rect 27433 2972 27445 2975
rect 27304 2944 27445 2972
rect 27304 2932 27310 2944
rect 27433 2941 27445 2944
rect 27479 2941 27491 2975
rect 32306 2972 32312 2984
rect 32267 2944 32312 2972
rect 27433 2935 27491 2941
rect 32306 2932 32312 2944
rect 32364 2932 32370 2984
rect 32398 2932 32404 2984
rect 32456 2972 32462 2984
rect 32585 2975 32643 2981
rect 32585 2972 32597 2975
rect 32456 2944 32597 2972
rect 32456 2932 32462 2944
rect 32585 2941 32597 2944
rect 32631 2941 32643 2975
rect 39298 2972 39304 2984
rect 39259 2944 39304 2972
rect 32585 2935 32643 2941
rect 39298 2932 39304 2944
rect 39356 2932 39362 2984
rect 5224 2876 8524 2904
rect 5224 2864 5230 2876
rect 13538 2864 13544 2916
rect 13596 2864 13602 2916
rect 38654 2904 38660 2916
rect 16546 2876 38660 2904
rect 6546 2796 6552 2848
rect 6604 2836 6610 2848
rect 6641 2839 6699 2845
rect 6641 2836 6653 2839
rect 6604 2808 6653 2836
rect 6604 2796 6610 2808
rect 6641 2805 6653 2808
rect 6687 2805 6699 2839
rect 6641 2799 6699 2805
rect 7377 2839 7435 2845
rect 7377 2805 7389 2839
rect 7423 2836 7435 2839
rect 8938 2836 8944 2848
rect 7423 2808 8944 2836
rect 7423 2805 7435 2808
rect 7377 2799 7435 2805
rect 8938 2796 8944 2808
rect 8996 2796 9002 2848
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 16546 2836 16574 2876
rect 38654 2864 38660 2876
rect 38712 2864 38718 2916
rect 9548 2808 16574 2836
rect 9548 2796 9554 2808
rect 18782 2796 18788 2848
rect 18840 2836 18846 2848
rect 39960 2836 39988 3012
rect 40770 3000 40776 3012
rect 40828 3040 40834 3052
rect 41693 3043 41751 3049
rect 41693 3040 41705 3043
rect 40828 3012 41705 3040
rect 40828 3000 40834 3012
rect 41693 3009 41705 3012
rect 41739 3009 41751 3043
rect 44726 3040 44732 3052
rect 44687 3012 44732 3040
rect 41693 3003 41751 3009
rect 44726 3000 44732 3012
rect 44784 3000 44790 3052
rect 47596 3049 47624 3080
rect 47581 3043 47639 3049
rect 47581 3009 47593 3043
rect 47627 3009 47639 3043
rect 47581 3003 47639 3009
rect 41049 2975 41107 2981
rect 41049 2941 41061 2975
rect 41095 2972 41107 2975
rect 42429 2975 42487 2981
rect 42429 2972 42441 2975
rect 41095 2944 42441 2972
rect 41095 2941 41107 2944
rect 41049 2935 41107 2941
rect 42429 2941 42441 2944
rect 42475 2941 42487 2975
rect 42429 2935 42487 2941
rect 42889 2975 42947 2981
rect 42889 2941 42901 2975
rect 42935 2941 42947 2975
rect 42889 2935 42947 2941
rect 41230 2864 41236 2916
rect 41288 2904 41294 2916
rect 42904 2904 42932 2935
rect 43622 2932 43628 2984
rect 43680 2972 43686 2984
rect 44913 2975 44971 2981
rect 44913 2972 44925 2975
rect 43680 2944 44925 2972
rect 43680 2932 43686 2944
rect 44913 2941 44925 2944
rect 44959 2941 44971 2975
rect 46566 2972 46572 2984
rect 46527 2944 46572 2972
rect 44913 2935 44971 2941
rect 46566 2932 46572 2944
rect 46624 2932 46630 2984
rect 41288 2876 42932 2904
rect 41288 2864 41294 2876
rect 43346 2864 43352 2916
rect 43404 2904 43410 2916
rect 45738 2904 45744 2916
rect 43404 2876 45744 2904
rect 43404 2864 43410 2876
rect 45738 2864 45744 2876
rect 45796 2864 45802 2916
rect 18840 2808 39988 2836
rect 41785 2839 41843 2845
rect 18840 2796 18846 2808
rect 41785 2805 41797 2839
rect 41831 2836 41843 2839
rect 42610 2836 42616 2848
rect 41831 2808 42616 2836
rect 41831 2805 41843 2808
rect 41785 2799 41843 2805
rect 42610 2796 42616 2808
rect 42668 2796 42674 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 1394 2592 1400 2644
rect 1452 2632 1458 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 1452 2604 2421 2632
rect 1452 2592 1458 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2409 2595 2467 2601
rect 19426 2592 19432 2644
rect 19484 2632 19490 2644
rect 19889 2635 19947 2641
rect 19889 2632 19901 2635
rect 19484 2604 19901 2632
rect 19484 2592 19490 2604
rect 19889 2601 19901 2604
rect 19935 2601 19947 2635
rect 19889 2595 19947 2601
rect 47486 2592 47492 2644
rect 47544 2632 47550 2644
rect 47765 2635 47823 2641
rect 47765 2632 47777 2635
rect 47544 2604 47777 2632
rect 47544 2592 47550 2604
rect 47765 2601 47777 2604
rect 47811 2601 47823 2635
rect 47765 2595 47823 2601
rect 1765 2567 1823 2573
rect 1765 2533 1777 2567
rect 1811 2564 1823 2567
rect 3786 2564 3792 2576
rect 1811 2536 3792 2564
rect 1811 2533 1823 2536
rect 1765 2527 1823 2533
rect 3786 2524 3792 2536
rect 3844 2524 3850 2576
rect 4522 2524 4528 2576
rect 4580 2564 4586 2576
rect 4580 2536 6868 2564
rect 4580 2524 4586 2536
rect 3326 2456 3332 2508
rect 3384 2496 3390 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 3384 2468 4261 2496
rect 3384 2456 3390 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 5868 2468 6377 2496
rect 5868 2456 5874 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6365 2459 6423 2465
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6840 2505 6868 2536
rect 7742 2524 7748 2576
rect 7800 2564 7806 2576
rect 27798 2564 27804 2576
rect 7800 2536 9444 2564
rect 7800 2524 7806 2536
rect 6825 2499 6883 2505
rect 6825 2465 6837 2499
rect 6871 2465 6883 2499
rect 8938 2496 8944 2508
rect 8899 2468 8944 2496
rect 6825 2459 6883 2465
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 9122 2496 9128 2508
rect 9083 2468 9128 2496
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 9416 2505 9444 2536
rect 27172 2536 27804 2564
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 27172 2505 27200 2536
rect 27798 2524 27804 2536
rect 27856 2524 27862 2576
rect 45830 2564 45836 2576
rect 45020 2536 45836 2564
rect 24673 2499 24731 2505
rect 24673 2496 24685 2499
rect 24268 2468 24685 2496
rect 24268 2456 24274 2468
rect 24673 2465 24685 2468
rect 24719 2465 24731 2499
rect 24673 2459 24731 2465
rect 27157 2499 27215 2505
rect 27157 2465 27169 2499
rect 27203 2465 27215 2499
rect 27157 2459 27215 2465
rect 27341 2499 27399 2505
rect 27341 2465 27353 2499
rect 27387 2496 27399 2499
rect 28350 2496 28356 2508
rect 27387 2468 28356 2496
rect 27387 2465 27399 2468
rect 27341 2459 27399 2465
rect 28350 2456 28356 2468
rect 28408 2456 28414 2508
rect 28537 2499 28595 2505
rect 28537 2465 28549 2499
rect 28583 2465 28595 2499
rect 28537 2459 28595 2465
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3283 2400 3801 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 23900 2400 24409 2428
rect 23900 2388 23906 2400
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 3973 2363 4031 2369
rect 3973 2329 3985 2363
rect 4019 2360 4031 2363
rect 4982 2360 4988 2372
rect 4019 2332 4988 2360
rect 4019 2329 4031 2332
rect 3973 2323 4031 2329
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 27706 2320 27712 2372
rect 27764 2360 27770 2372
rect 28552 2360 28580 2459
rect 42334 2456 42340 2508
rect 42392 2496 42398 2508
rect 42429 2499 42487 2505
rect 42429 2496 42441 2499
rect 42392 2468 42441 2496
rect 42392 2456 42398 2468
rect 42429 2465 42441 2468
rect 42475 2465 42487 2499
rect 42610 2496 42616 2508
rect 42571 2468 42616 2496
rect 42429 2459 42487 2465
rect 42610 2456 42616 2468
rect 42668 2456 42674 2508
rect 45020 2505 45048 2536
rect 45830 2524 45836 2536
rect 45888 2524 45894 2576
rect 45005 2499 45063 2505
rect 45005 2465 45017 2499
rect 45051 2465 45063 2499
rect 45186 2496 45192 2508
rect 45147 2468 45192 2496
rect 45005 2459 45063 2465
rect 45186 2456 45192 2468
rect 45244 2456 45250 2508
rect 45278 2456 45284 2508
rect 45336 2496 45342 2508
rect 45557 2499 45615 2505
rect 45557 2496 45569 2499
rect 45336 2468 45569 2496
rect 45336 2456 45342 2468
rect 45557 2465 45569 2468
rect 45603 2465 45615 2499
rect 45557 2459 45615 2465
rect 27764 2332 28580 2360
rect 44269 2363 44327 2369
rect 27764 2320 27770 2332
rect 44269 2329 44281 2363
rect 44315 2360 44327 2363
rect 48958 2360 48964 2372
rect 44315 2332 48964 2360
rect 44315 2329 44327 2332
rect 44269 2323 44327 2329
rect 48958 2320 48964 2332
rect 49016 2320 49022 2372
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
<< via1 >>
rect 38660 47404 38712 47456
rect 39948 47404 40000 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 2964 47132 3016 47184
rect 27620 47132 27672 47184
rect 45192 47132 45244 47184
rect 20 47064 72 47116
rect 2688 46996 2740 47048
rect 11520 47064 11572 47116
rect 28816 47064 28868 47116
rect 46848 47064 46900 47116
rect 4252 47039 4304 47048
rect 4252 47005 4261 47039
rect 4261 47005 4295 47039
rect 4295 47005 4304 47039
rect 4252 46996 4304 47005
rect 5540 47039 5592 47048
rect 5540 47005 5549 47039
rect 5549 47005 5583 47039
rect 5583 47005 5592 47039
rect 5540 46996 5592 47005
rect 8392 46996 8444 47048
rect 12716 47039 12768 47048
rect 12716 47005 12725 47039
rect 12725 47005 12759 47039
rect 12759 47005 12768 47039
rect 12716 46996 12768 47005
rect 13176 46996 13228 47048
rect 14188 46996 14240 47048
rect 15660 47039 15712 47048
rect 15660 47005 15669 47039
rect 15669 47005 15703 47039
rect 15703 47005 15712 47039
rect 15660 46996 15712 47005
rect 24860 47039 24912 47048
rect 24860 47005 24869 47039
rect 24869 47005 24903 47039
rect 24903 47005 24912 47039
rect 24860 46996 24912 47005
rect 25504 47039 25556 47048
rect 25504 47005 25513 47039
rect 25513 47005 25547 47039
rect 25547 47005 25556 47039
rect 25504 46996 25556 47005
rect 26424 47039 26476 47048
rect 26424 47005 26433 47039
rect 26433 47005 26467 47039
rect 26467 47005 26476 47039
rect 26424 46996 26476 47005
rect 27988 47039 28040 47048
rect 27988 47005 27997 47039
rect 27997 47005 28031 47039
rect 28031 47005 28040 47039
rect 27988 46996 28040 47005
rect 29736 46996 29788 47048
rect 32772 46996 32824 47048
rect 37280 46996 37332 47048
rect 46388 47039 46440 47048
rect 46388 47005 46397 47039
rect 46397 47005 46431 47039
rect 46431 47005 46440 47039
rect 46388 46996 46440 47005
rect 47124 46996 47176 47048
rect 2872 46971 2924 46980
rect 2872 46937 2881 46971
rect 2881 46937 2915 46971
rect 2915 46937 2924 46971
rect 2872 46928 2924 46937
rect 46572 46928 46624 46980
rect 8944 46903 8996 46912
rect 8944 46869 8953 46903
rect 8953 46869 8987 46903
rect 8987 46869 8996 46903
rect 8944 46860 8996 46869
rect 40592 46860 40644 46912
rect 41420 46860 41472 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 2596 46656 2648 46708
rect 3056 46656 3108 46708
rect 3884 46588 3936 46640
rect 4252 46588 4304 46640
rect 12716 46588 12768 46640
rect 14188 46563 14240 46572
rect 14188 46529 14197 46563
rect 14197 46529 14231 46563
rect 14231 46529 14240 46563
rect 14188 46520 14240 46529
rect 25504 46588 25556 46640
rect 26424 46520 26476 46572
rect 29736 46563 29788 46572
rect 29736 46529 29745 46563
rect 29745 46529 29779 46563
rect 29779 46529 29788 46563
rect 29736 46520 29788 46529
rect 32772 46563 32824 46572
rect 32772 46529 32781 46563
rect 32781 46529 32815 46563
rect 32815 46529 32824 46563
rect 32772 46520 32824 46529
rect 35808 46563 35860 46572
rect 35808 46529 35817 46563
rect 35817 46529 35851 46563
rect 35851 46529 35860 46563
rect 35808 46520 35860 46529
rect 37280 46563 37332 46572
rect 37280 46529 37289 46563
rect 37289 46529 37323 46563
rect 37323 46529 37332 46563
rect 37280 46520 37332 46529
rect 46388 46588 46440 46640
rect 47216 46520 47268 46572
rect 2136 46495 2188 46504
rect 2136 46461 2145 46495
rect 2145 46461 2179 46495
rect 2179 46461 2188 46495
rect 2136 46452 2188 46461
rect 4620 46495 4672 46504
rect 1768 46384 1820 46436
rect 4068 46384 4120 46436
rect 4620 46461 4629 46495
rect 4629 46461 4663 46495
rect 4663 46461 4672 46495
rect 4620 46452 4672 46461
rect 12624 46452 12676 46504
rect 12900 46495 12952 46504
rect 12900 46461 12909 46495
rect 12909 46461 12943 46495
rect 12943 46461 12952 46495
rect 12900 46452 12952 46461
rect 14464 46452 14516 46504
rect 14832 46495 14884 46504
rect 14832 46461 14841 46495
rect 14841 46461 14875 46495
rect 14875 46461 14884 46495
rect 14832 46452 14884 46461
rect 22284 46495 22336 46504
rect 22284 46461 22293 46495
rect 22293 46461 22327 46495
rect 22327 46461 22336 46495
rect 22284 46452 22336 46461
rect 22928 46452 22980 46504
rect 23204 46495 23256 46504
rect 23204 46461 23213 46495
rect 23213 46461 23247 46495
rect 23247 46461 23256 46495
rect 23204 46452 23256 46461
rect 25320 46452 25372 46504
rect 25780 46495 25832 46504
rect 25780 46461 25789 46495
rect 25789 46461 25823 46495
rect 25823 46461 25832 46495
rect 25780 46452 25832 46461
rect 26240 46452 26292 46504
rect 29920 46495 29972 46504
rect 9588 46384 9640 46436
rect 17224 46384 17276 46436
rect 27068 46384 27120 46436
rect 29920 46461 29929 46495
rect 29929 46461 29963 46495
rect 29963 46461 29972 46495
rect 29920 46452 29972 46461
rect 30288 46452 30340 46504
rect 32956 46495 33008 46504
rect 32956 46461 32965 46495
rect 32965 46461 32999 46495
rect 32999 46461 33008 46495
rect 32956 46452 33008 46461
rect 33508 46495 33560 46504
rect 33508 46461 33517 46495
rect 33517 46461 33551 46495
rect 33551 46461 33560 46495
rect 33508 46452 33560 46461
rect 37464 46495 37516 46504
rect 37464 46461 37473 46495
rect 37473 46461 37507 46495
rect 37507 46461 37516 46495
rect 37464 46452 37516 46461
rect 35716 46384 35768 46436
rect 36728 46384 36780 46436
rect 46572 46452 46624 46504
rect 46756 46495 46808 46504
rect 46756 46461 46765 46495
rect 46765 46461 46799 46495
rect 46799 46461 46808 46495
rect 46756 46452 46808 46461
rect 10876 46316 10928 46368
rect 35900 46359 35952 46368
rect 35900 46325 35909 46359
rect 35909 46325 35943 46359
rect 35943 46325 35952 46359
rect 35900 46316 35952 46325
rect 41604 46316 41656 46368
rect 45652 46316 45704 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 4068 46112 4120 46164
rect 14464 46155 14516 46164
rect 14464 46121 14473 46155
rect 14473 46121 14507 46155
rect 14507 46121 14516 46155
rect 14464 46112 14516 46121
rect 22284 46112 22336 46164
rect 32956 46112 33008 46164
rect 10968 46044 11020 46096
rect 15476 46044 15528 46096
rect 2780 46019 2832 46028
rect 2780 45985 2789 46019
rect 2789 45985 2823 46019
rect 2823 45985 2832 46019
rect 2780 45976 2832 45985
rect 5540 45976 5592 46028
rect 5816 46019 5868 46028
rect 5816 45985 5825 46019
rect 5825 45985 5859 46019
rect 5859 45985 5868 46019
rect 5816 45976 5868 45985
rect 9588 46019 9640 46028
rect 9588 45985 9597 46019
rect 9597 45985 9631 46019
rect 9631 45985 9640 46019
rect 9588 45976 9640 45985
rect 10876 46019 10928 46028
rect 10876 45985 10885 46019
rect 10885 45985 10919 46019
rect 10919 45985 10928 46019
rect 10876 45976 10928 45985
rect 15660 45976 15712 46028
rect 17224 45976 17276 46028
rect 47216 46112 47268 46164
rect 36084 45976 36136 46028
rect 41604 46019 41656 46028
rect 41604 45985 41613 46019
rect 41613 45985 41647 46019
rect 41647 45985 41656 46019
rect 41604 45976 41656 45985
rect 42064 46019 42116 46028
rect 42064 45985 42073 46019
rect 42073 45985 42107 46019
rect 42107 45985 42116 46019
rect 42064 45976 42116 45985
rect 48320 45976 48372 46028
rect 1400 45951 1452 45960
rect 1400 45917 1409 45951
rect 1409 45917 1443 45951
rect 1443 45917 1452 45951
rect 1400 45908 1452 45917
rect 9220 45951 9272 45960
rect 3148 45840 3200 45892
rect 9220 45917 9229 45951
rect 9229 45917 9263 45951
rect 9263 45917 9272 45951
rect 9220 45908 9272 45917
rect 12532 45908 12584 45960
rect 24676 45951 24728 45960
rect 5540 45840 5592 45892
rect 11612 45840 11664 45892
rect 24676 45917 24685 45951
rect 24685 45917 24719 45951
rect 24719 45917 24728 45951
rect 24676 45908 24728 45917
rect 26976 45951 27028 45960
rect 26976 45917 26985 45951
rect 26985 45917 27019 45951
rect 27019 45917 27028 45951
rect 26976 45908 27028 45917
rect 28816 45951 28868 45960
rect 28816 45917 28825 45951
rect 28825 45917 28859 45951
rect 28859 45917 28868 45951
rect 28816 45908 28868 45917
rect 29736 45951 29788 45960
rect 29736 45917 29745 45951
rect 29745 45917 29779 45951
rect 29779 45917 29788 45951
rect 29736 45908 29788 45917
rect 32772 45951 32824 45960
rect 32772 45917 32781 45951
rect 32781 45917 32815 45951
rect 32815 45917 32824 45951
rect 32772 45908 32824 45917
rect 35716 45951 35768 45960
rect 35716 45917 35725 45951
rect 35725 45917 35759 45951
rect 35759 45917 35768 45951
rect 35716 45908 35768 45917
rect 38108 45908 38160 45960
rect 15568 45883 15620 45892
rect 15568 45849 15577 45883
rect 15577 45849 15611 45883
rect 15611 45849 15620 45883
rect 15568 45840 15620 45849
rect 24860 45883 24912 45892
rect 24860 45849 24869 45883
rect 24869 45849 24903 45883
rect 24903 45849 24912 45883
rect 24860 45840 24912 45849
rect 25136 45840 25188 45892
rect 27160 45883 27212 45892
rect 27160 45849 27169 45883
rect 27169 45849 27203 45883
rect 27203 45849 27212 45883
rect 27160 45840 27212 45849
rect 35900 45883 35952 45892
rect 35900 45849 35909 45883
rect 35909 45849 35943 45883
rect 35943 45849 35952 45883
rect 41788 45883 41840 45892
rect 35900 45840 35952 45849
rect 41788 45849 41797 45883
rect 41797 45849 41831 45883
rect 41831 45849 41840 45883
rect 41788 45840 41840 45849
rect 47676 45840 47728 45892
rect 4068 45772 4120 45824
rect 10784 45772 10836 45824
rect 13360 45772 13412 45824
rect 14372 45772 14424 45824
rect 35808 45772 35860 45824
rect 40684 45772 40736 45824
rect 47124 45772 47176 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 11612 45611 11664 45620
rect 11612 45577 11621 45611
rect 11621 45577 11655 45611
rect 11655 45577 11664 45611
rect 11612 45568 11664 45577
rect 1676 45543 1728 45552
rect 1676 45509 1685 45543
rect 1685 45509 1719 45543
rect 1719 45509 1728 45543
rect 1676 45500 1728 45509
rect 2872 45500 2924 45552
rect 5540 45543 5592 45552
rect 5540 45509 5549 45543
rect 5549 45509 5583 45543
rect 5583 45509 5592 45543
rect 5540 45500 5592 45509
rect 5448 45475 5500 45484
rect 5448 45441 5457 45475
rect 5457 45441 5491 45475
rect 5491 45441 5500 45475
rect 9588 45500 9640 45552
rect 12624 45543 12676 45552
rect 12624 45509 12633 45543
rect 12633 45509 12667 45543
rect 12667 45509 12676 45543
rect 12624 45500 12676 45509
rect 13360 45543 13412 45552
rect 8392 45475 8444 45484
rect 5448 45432 5500 45441
rect 8392 45441 8401 45475
rect 8401 45441 8435 45475
rect 8435 45441 8444 45475
rect 8392 45432 8444 45441
rect 9220 45432 9272 45484
rect 11520 45475 11572 45484
rect 11520 45441 11529 45475
rect 11529 45441 11563 45475
rect 11563 45441 11572 45475
rect 11520 45432 11572 45441
rect 12532 45475 12584 45484
rect 12532 45441 12541 45475
rect 12541 45441 12575 45475
rect 12575 45441 12584 45475
rect 12532 45432 12584 45441
rect 2964 45364 3016 45416
rect 3056 45407 3108 45416
rect 3056 45373 3065 45407
rect 3065 45373 3099 45407
rect 3099 45373 3108 45407
rect 9404 45407 9456 45416
rect 3056 45364 3108 45373
rect 9404 45373 9413 45407
rect 9413 45373 9447 45407
rect 9447 45373 9456 45407
rect 9404 45364 9456 45373
rect 10784 45364 10836 45416
rect 13360 45509 13369 45543
rect 13369 45509 13403 45543
rect 13403 45509 13412 45543
rect 13360 45500 13412 45509
rect 15568 45568 15620 45620
rect 22928 45611 22980 45620
rect 22928 45577 22937 45611
rect 22937 45577 22971 45611
rect 22971 45577 22980 45611
rect 22928 45568 22980 45577
rect 32772 45568 32824 45620
rect 40684 45568 40736 45620
rect 18512 45500 18564 45552
rect 24860 45500 24912 45552
rect 25320 45543 25372 45552
rect 25320 45509 25329 45543
rect 25329 45509 25363 45543
rect 25363 45509 25372 45543
rect 25320 45500 25372 45509
rect 13176 45475 13228 45484
rect 13176 45441 13185 45475
rect 13185 45441 13219 45475
rect 13219 45441 13228 45475
rect 13176 45432 13228 45441
rect 15568 45475 15620 45484
rect 15568 45441 15577 45475
rect 15577 45441 15611 45475
rect 15611 45441 15620 45475
rect 22836 45475 22888 45484
rect 15568 45432 15620 45441
rect 14280 45407 14332 45416
rect 8392 45296 8444 45348
rect 14280 45373 14289 45407
rect 14289 45373 14323 45407
rect 14323 45373 14332 45407
rect 14280 45364 14332 45373
rect 22836 45441 22845 45475
rect 22845 45441 22879 45475
rect 22879 45441 22888 45475
rect 22836 45432 22888 45441
rect 24492 45432 24544 45484
rect 26240 45432 26292 45484
rect 26976 45432 27028 45484
rect 26056 45296 26108 45348
rect 29736 45500 29788 45552
rect 39948 45543 40000 45552
rect 39948 45509 39957 45543
rect 39957 45509 39991 45543
rect 39991 45509 40000 45543
rect 39948 45500 40000 45509
rect 45652 45500 45704 45552
rect 47676 45543 47728 45552
rect 47676 45509 47685 45543
rect 47685 45509 47719 45543
rect 47719 45509 47728 45543
rect 47676 45500 47728 45509
rect 36084 45432 36136 45484
rect 38108 45475 38160 45484
rect 38108 45441 38117 45475
rect 38117 45441 38151 45475
rect 38151 45441 38160 45475
rect 38108 45432 38160 45441
rect 45192 45475 45244 45484
rect 45192 45441 45201 45475
rect 45201 45441 45235 45475
rect 45235 45441 45244 45475
rect 45192 45432 45244 45441
rect 47308 45432 47360 45484
rect 27436 45364 27488 45416
rect 30288 45407 30340 45416
rect 30288 45373 30297 45407
rect 30297 45373 30331 45407
rect 30331 45373 30340 45407
rect 30288 45364 30340 45373
rect 38016 45364 38068 45416
rect 38292 45407 38344 45416
rect 38292 45373 38301 45407
rect 38301 45373 38335 45407
rect 38335 45373 38344 45407
rect 38292 45364 38344 45373
rect 46848 45407 46900 45416
rect 46848 45373 46857 45407
rect 46857 45373 46891 45407
rect 46891 45373 46900 45407
rect 46848 45364 46900 45373
rect 37464 45296 37516 45348
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 1400 45024 1452 45076
rect 3148 45067 3200 45076
rect 3148 45033 3157 45067
rect 3157 45033 3191 45067
rect 3191 45033 3200 45067
rect 3148 45024 3200 45033
rect 3884 45067 3936 45076
rect 3884 45033 3893 45067
rect 3893 45033 3927 45067
rect 3927 45033 3936 45067
rect 3884 45024 3936 45033
rect 27160 45024 27212 45076
rect 27436 45067 27488 45076
rect 27436 45033 27445 45067
rect 27445 45033 27479 45067
rect 27479 45033 27488 45067
rect 27436 45024 27488 45033
rect 29920 45024 29972 45076
rect 38292 45024 38344 45076
rect 41788 45067 41840 45076
rect 41788 45033 41797 45067
rect 41797 45033 41831 45067
rect 41831 45033 41840 45067
rect 41788 45024 41840 45033
rect 1768 44956 1820 45008
rect 9404 44956 9456 45008
rect 3056 44863 3108 44872
rect 3056 44829 3065 44863
rect 3065 44829 3099 44863
rect 3099 44829 3108 44863
rect 3056 44820 3108 44829
rect 8208 44888 8260 44940
rect 14372 44888 14424 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 9220 44863 9272 44872
rect 9220 44829 9229 44863
rect 9229 44829 9263 44863
rect 9263 44829 9272 44863
rect 9220 44820 9272 44829
rect 26700 44863 26752 44872
rect 26700 44829 26709 44863
rect 26709 44829 26743 44863
rect 26743 44829 26752 44863
rect 26700 44820 26752 44829
rect 29920 44863 29972 44872
rect 29920 44829 29929 44863
rect 29929 44829 29963 44863
rect 29963 44829 29972 44863
rect 29920 44820 29972 44829
rect 38292 44820 38344 44872
rect 41972 44820 42024 44872
rect 9588 44795 9640 44804
rect 9588 44761 9597 44795
rect 9597 44761 9631 44795
rect 9631 44761 9640 44795
rect 9588 44752 9640 44761
rect 22836 44752 22888 44804
rect 46480 44795 46532 44804
rect 46480 44761 46489 44795
rect 46489 44761 46523 44795
rect 46523 44761 46532 44795
rect 46480 44752 46532 44761
rect 38292 44684 38344 44736
rect 47584 44684 47636 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 3056 44480 3108 44532
rect 15568 44480 15620 44532
rect 46480 44480 46532 44532
rect 29920 44412 29972 44464
rect 9220 44344 9272 44396
rect 38016 44344 38068 44396
rect 47860 44344 47912 44396
rect 9036 44276 9088 44328
rect 32772 44276 32824 44328
rect 45376 44208 45428 44260
rect 45192 44140 45244 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 48044 43843 48096 43852
rect 48044 43809 48053 43843
rect 48053 43809 48087 43843
rect 48087 43809 48096 43843
rect 48044 43800 48096 43809
rect 2136 43732 2188 43784
rect 40040 43732 40092 43784
rect 46020 43732 46072 43784
rect 46572 43664 46624 43716
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 46572 43435 46624 43444
rect 46572 43401 46581 43435
rect 46581 43401 46615 43435
rect 46615 43401 46624 43435
rect 46572 43392 46624 43401
rect 3976 43367 4028 43376
rect 3976 43333 3985 43367
rect 3985 43333 4019 43367
rect 4019 43333 4028 43367
rect 3976 43324 4028 43333
rect 2136 43299 2188 43308
rect 2136 43265 2145 43299
rect 2145 43265 2179 43299
rect 2179 43265 2188 43299
rect 2136 43256 2188 43265
rect 40040 43299 40092 43308
rect 40040 43265 40049 43299
rect 40049 43265 40083 43299
rect 40083 43265 40092 43299
rect 40040 43256 40092 43265
rect 46020 43299 46072 43308
rect 46020 43265 46029 43299
rect 46029 43265 46063 43299
rect 46063 43265 46072 43299
rect 46020 43256 46072 43265
rect 46480 43299 46532 43308
rect 46480 43265 46489 43299
rect 46489 43265 46523 43299
rect 46523 43265 46532 43299
rect 46480 43256 46532 43265
rect 47584 43299 47636 43308
rect 47584 43265 47593 43299
rect 47593 43265 47627 43299
rect 47627 43265 47636 43299
rect 47584 43256 47636 43265
rect 3884 43188 3936 43240
rect 40224 43231 40276 43240
rect 40224 43197 40233 43231
rect 40233 43197 40267 43231
rect 40267 43197 40276 43231
rect 40224 43188 40276 43197
rect 41420 43231 41472 43240
rect 41420 43197 41429 43231
rect 41429 43197 41463 43231
rect 41463 43197 41472 43231
rect 41420 43188 41472 43197
rect 47676 43095 47728 43104
rect 47676 43061 47685 43095
rect 47685 43061 47719 43095
rect 47719 43061 47728 43095
rect 47676 43052 47728 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 3884 42755 3936 42764
rect 3884 42721 3893 42755
rect 3893 42721 3927 42755
rect 3927 42721 3936 42755
rect 3884 42712 3936 42721
rect 30656 42712 30708 42764
rect 47676 42712 47728 42764
rect 6368 42644 6420 42696
rect 9588 42644 9640 42696
rect 27620 42644 27672 42696
rect 8944 42576 8996 42628
rect 33784 42644 33836 42696
rect 45744 42644 45796 42696
rect 48136 42619 48188 42628
rect 48136 42585 48145 42619
rect 48145 42585 48179 42619
rect 48179 42585 48188 42619
rect 48136 42576 48188 42585
rect 27160 42508 27212 42560
rect 28540 42508 28592 42560
rect 33508 42551 33560 42560
rect 33508 42517 33517 42551
rect 33517 42517 33551 42551
rect 33551 42517 33560 42551
rect 33508 42508 33560 42517
rect 45284 42508 45336 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 40224 42304 40276 42356
rect 33508 42236 33560 42288
rect 27160 42211 27212 42220
rect 27160 42177 27169 42211
rect 27169 42177 27203 42211
rect 27203 42177 27212 42211
rect 27160 42168 27212 42177
rect 28540 42211 28592 42220
rect 28540 42177 28549 42211
rect 28549 42177 28583 42211
rect 28583 42177 28592 42211
rect 28540 42168 28592 42177
rect 31392 42211 31444 42220
rect 31392 42177 31401 42211
rect 31401 42177 31435 42211
rect 31435 42177 31444 42211
rect 31392 42168 31444 42177
rect 32680 42211 32732 42220
rect 32680 42177 32689 42211
rect 32689 42177 32723 42211
rect 32723 42177 32732 42211
rect 32680 42168 32732 42177
rect 45376 42279 45428 42288
rect 45376 42245 45385 42279
rect 45385 42245 45419 42279
rect 45419 42245 45428 42279
rect 45376 42236 45428 42245
rect 33140 42143 33192 42152
rect 33140 42109 33149 42143
rect 33149 42109 33183 42143
rect 33183 42109 33192 42143
rect 33140 42100 33192 42109
rect 26976 42007 27028 42016
rect 26976 41973 26985 42007
rect 26985 41973 27019 42007
rect 27019 41973 27028 42007
rect 26976 41964 27028 41973
rect 29644 41964 29696 42016
rect 31208 42007 31260 42016
rect 31208 41973 31217 42007
rect 31217 41973 31251 42007
rect 31251 41973 31260 42007
rect 31208 41964 31260 41973
rect 32496 42007 32548 42016
rect 32496 41973 32505 42007
rect 32505 41973 32539 42007
rect 32539 41973 32548 42007
rect 32496 41964 32548 41973
rect 34520 42007 34572 42016
rect 34520 41973 34529 42007
rect 34529 41973 34563 42007
rect 34563 41973 34572 42007
rect 36728 42100 36780 42152
rect 38200 42168 38252 42220
rect 41144 42168 41196 42220
rect 41604 42211 41656 42220
rect 41604 42177 41613 42211
rect 41613 42177 41647 42211
rect 41647 42177 41656 42211
rect 41604 42168 41656 42177
rect 42524 42211 42576 42220
rect 42524 42177 42533 42211
rect 42533 42177 42567 42211
rect 42567 42177 42576 42211
rect 42524 42168 42576 42177
rect 45192 42211 45244 42220
rect 45192 42177 45201 42211
rect 45201 42177 45235 42211
rect 45235 42177 45244 42211
rect 45192 42168 45244 42177
rect 46848 42143 46900 42152
rect 46848 42109 46857 42143
rect 46857 42109 46891 42143
rect 46891 42109 46900 42143
rect 46848 42100 46900 42109
rect 40224 42032 40276 42084
rect 34520 41964 34572 41973
rect 35348 41964 35400 42016
rect 35808 42007 35860 42016
rect 35808 41973 35817 42007
rect 35817 41973 35851 42007
rect 35851 41973 35860 42007
rect 35808 41964 35860 41973
rect 36452 42007 36504 42016
rect 36452 41973 36461 42007
rect 36461 41973 36495 42007
rect 36495 41973 36504 42007
rect 36452 41964 36504 41973
rect 41880 42007 41932 42016
rect 41880 41973 41889 42007
rect 41889 41973 41923 42007
rect 41923 41973 41932 42007
rect 41880 41964 41932 41973
rect 43260 42007 43312 42016
rect 43260 41973 43269 42007
rect 43269 41973 43303 42007
rect 43303 41973 43312 42007
rect 43260 41964 43312 41973
rect 46296 41964 46348 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 32680 41760 32732 41812
rect 36728 41760 36780 41812
rect 42524 41803 42576 41812
rect 42524 41769 42533 41803
rect 42533 41769 42567 41803
rect 42567 41769 42576 41803
rect 42524 41760 42576 41769
rect 29552 41599 29604 41608
rect 29552 41565 29561 41599
rect 29561 41565 29595 41599
rect 29595 41565 29604 41599
rect 29552 41556 29604 41565
rect 29644 41556 29696 41608
rect 33140 41556 33192 41608
rect 26976 41488 27028 41540
rect 31208 41488 31260 41540
rect 33600 41556 33652 41608
rect 35808 41556 35860 41608
rect 37648 41556 37700 41608
rect 27896 41463 27948 41472
rect 27896 41429 27905 41463
rect 27905 41429 27939 41463
rect 27939 41429 27948 41463
rect 27896 41420 27948 41429
rect 30932 41463 30984 41472
rect 30932 41429 30941 41463
rect 30941 41429 30975 41463
rect 30975 41429 30984 41463
rect 30932 41420 30984 41429
rect 34612 41488 34664 41540
rect 36452 41488 36504 41540
rect 39396 41556 39448 41608
rect 40224 41624 40276 41676
rect 46296 41667 46348 41676
rect 46296 41633 46305 41667
rect 46305 41633 46339 41667
rect 46339 41633 46348 41667
rect 46296 41624 46348 41633
rect 40132 41556 40184 41608
rect 43996 41556 44048 41608
rect 45100 41599 45152 41608
rect 45100 41565 45109 41599
rect 45109 41565 45143 41599
rect 45143 41565 45152 41599
rect 45100 41556 45152 41565
rect 45284 41599 45336 41608
rect 45284 41565 45293 41599
rect 45293 41565 45327 41599
rect 45327 41565 45336 41599
rect 45284 41556 45336 41565
rect 41696 41488 41748 41540
rect 43260 41531 43312 41540
rect 43260 41497 43294 41531
rect 43294 41497 43312 41531
rect 43260 41488 43312 41497
rect 46940 41488 46992 41540
rect 48228 41488 48280 41540
rect 38108 41420 38160 41472
rect 40040 41420 40092 41472
rect 43812 41420 43864 41472
rect 46020 41420 46072 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 31392 41216 31444 41268
rect 34428 41259 34480 41268
rect 32496 41148 32548 41200
rect 16948 41123 17000 41132
rect 16948 41089 16957 41123
rect 16957 41089 16991 41123
rect 16991 41089 17000 41123
rect 16948 41080 17000 41089
rect 8852 41055 8904 41064
rect 8852 41021 8861 41055
rect 8861 41021 8895 41055
rect 8895 41021 8904 41055
rect 8852 41012 8904 41021
rect 25964 41055 26016 41064
rect 3424 40944 3476 40996
rect 25964 41021 25973 41055
rect 25973 41021 26007 41055
rect 26007 41021 26016 41055
rect 25964 41012 26016 41021
rect 27068 41080 27120 41132
rect 29000 41080 29052 41132
rect 30012 41080 30064 41132
rect 34428 41225 34437 41259
rect 34437 41225 34471 41259
rect 34471 41225 34480 41259
rect 34428 41216 34480 41225
rect 39396 41259 39448 41268
rect 39396 41225 39405 41259
rect 39405 41225 39439 41259
rect 39439 41225 39448 41259
rect 39396 41216 39448 41225
rect 40040 41216 40092 41268
rect 41696 41259 41748 41268
rect 34520 41191 34572 41200
rect 34520 41157 34529 41191
rect 34529 41157 34563 41191
rect 34563 41157 34572 41191
rect 34520 41148 34572 41157
rect 34704 41148 34756 41200
rect 26608 41012 26660 41064
rect 30932 41012 30984 41064
rect 34796 41080 34848 41132
rect 37372 41148 37424 41200
rect 37648 41148 37700 41200
rect 41696 41225 41705 41259
rect 41705 41225 41739 41259
rect 41739 41225 41748 41259
rect 41696 41216 41748 41225
rect 42984 41216 43036 41268
rect 46940 41259 46992 41268
rect 46940 41225 46949 41259
rect 46949 41225 46983 41259
rect 46983 41225 46992 41259
rect 46940 41216 46992 41225
rect 37004 41080 37056 41132
rect 37556 41123 37608 41132
rect 37556 41089 37565 41123
rect 37565 41089 37599 41123
rect 37599 41089 37608 41123
rect 37556 41080 37608 41089
rect 35348 41055 35400 41064
rect 24584 40944 24636 40996
rect 25320 40919 25372 40928
rect 25320 40885 25329 40919
rect 25329 40885 25363 40919
rect 25363 40885 25372 40919
rect 25320 40876 25372 40885
rect 29368 40919 29420 40928
rect 29368 40885 29377 40919
rect 29377 40885 29411 40919
rect 29411 40885 29420 40919
rect 29368 40876 29420 40885
rect 35348 41021 35357 41055
rect 35357 41021 35391 41055
rect 35391 41021 35400 41055
rect 35348 41012 35400 41021
rect 42524 41148 42576 41200
rect 41880 41123 41932 41132
rect 41880 41089 41889 41123
rect 41889 41089 41923 41123
rect 41923 41089 41932 41123
rect 41880 41080 41932 41089
rect 33876 40944 33928 40996
rect 33140 40876 33192 40928
rect 33692 40876 33744 40928
rect 34428 40944 34480 40996
rect 34612 40876 34664 40928
rect 34796 40919 34848 40928
rect 34796 40885 34805 40919
rect 34805 40885 34839 40919
rect 34839 40885 34848 40919
rect 34796 40876 34848 40885
rect 35716 40919 35768 40928
rect 35716 40885 35725 40919
rect 35725 40885 35759 40919
rect 35759 40885 35768 40919
rect 35716 40876 35768 40885
rect 36544 40919 36596 40928
rect 36544 40885 36553 40919
rect 36553 40885 36587 40919
rect 36587 40885 36596 40919
rect 36544 40876 36596 40885
rect 36728 40919 36780 40928
rect 36728 40885 36737 40919
rect 36737 40885 36771 40919
rect 36771 40885 36780 40919
rect 36728 40876 36780 40885
rect 37464 40876 37516 40928
rect 41604 41012 41656 41064
rect 43812 41080 43864 41132
rect 43996 41123 44048 41132
rect 43996 41089 44005 41123
rect 44005 41089 44039 41123
rect 44039 41089 44048 41123
rect 43996 41080 44048 41089
rect 44088 41080 44140 41132
rect 46020 41123 46072 41132
rect 46020 41089 46029 41123
rect 46029 41089 46063 41123
rect 46063 41089 46072 41123
rect 46020 41080 46072 41089
rect 46664 41080 46716 41132
rect 40132 40876 40184 40928
rect 41236 40919 41288 40928
rect 41236 40885 41245 40919
rect 41245 40885 41279 40919
rect 41279 40885 41288 40919
rect 41236 40876 41288 40885
rect 42800 40876 42852 40928
rect 45836 40919 45888 40928
rect 45836 40885 45845 40919
rect 45845 40885 45879 40919
rect 45879 40885 45888 40919
rect 45836 40876 45888 40885
rect 46296 40876 46348 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 8852 40672 8904 40724
rect 25964 40672 26016 40724
rect 27896 40715 27948 40724
rect 27896 40681 27905 40715
rect 27905 40681 27939 40715
rect 27939 40681 27948 40715
rect 27896 40672 27948 40681
rect 29000 40715 29052 40724
rect 29000 40681 29009 40715
rect 29009 40681 29043 40715
rect 29043 40681 29052 40715
rect 29000 40672 29052 40681
rect 27252 40604 27304 40656
rect 32588 40672 32640 40724
rect 33784 40715 33836 40724
rect 33784 40681 33793 40715
rect 33793 40681 33827 40715
rect 33827 40681 33836 40715
rect 33784 40672 33836 40681
rect 37556 40672 37608 40724
rect 40224 40672 40276 40724
rect 41604 40715 41656 40724
rect 37648 40604 37700 40656
rect 41604 40681 41613 40715
rect 41613 40681 41647 40715
rect 41647 40681 41656 40715
rect 41604 40672 41656 40681
rect 2688 40536 2740 40588
rect 29552 40579 29604 40588
rect 29552 40545 29561 40579
rect 29561 40545 29595 40579
rect 29595 40545 29604 40579
rect 29552 40536 29604 40545
rect 24584 40511 24636 40520
rect 24584 40477 24593 40511
rect 24593 40477 24627 40511
rect 24627 40477 24636 40511
rect 24584 40468 24636 40477
rect 24860 40468 24912 40520
rect 25320 40511 25372 40520
rect 25320 40477 25354 40511
rect 25354 40477 25372 40511
rect 25320 40468 25372 40477
rect 23848 40400 23900 40452
rect 27068 40511 27120 40520
rect 27068 40477 27077 40511
rect 27077 40477 27111 40511
rect 27111 40477 27120 40511
rect 27896 40511 27948 40520
rect 27068 40468 27120 40477
rect 27896 40477 27905 40511
rect 27905 40477 27939 40511
rect 27939 40477 27948 40511
rect 27896 40468 27948 40477
rect 27988 40511 28040 40520
rect 27988 40477 27997 40511
rect 27997 40477 28031 40511
rect 28031 40477 28040 40511
rect 27988 40468 28040 40477
rect 27712 40443 27764 40452
rect 23480 40375 23532 40384
rect 23480 40341 23489 40375
rect 23489 40341 23523 40375
rect 23523 40341 23532 40375
rect 23480 40332 23532 40341
rect 24400 40375 24452 40384
rect 24400 40341 24409 40375
rect 24409 40341 24443 40375
rect 24443 40341 24452 40375
rect 24400 40332 24452 40341
rect 27712 40409 27721 40443
rect 27721 40409 27755 40443
rect 27755 40409 27764 40443
rect 27712 40400 27764 40409
rect 29184 40400 29236 40452
rect 29368 40468 29420 40520
rect 30012 40400 30064 40452
rect 33600 40511 33652 40520
rect 33600 40477 33609 40511
rect 33609 40477 33643 40511
rect 33643 40477 33652 40511
rect 36728 40536 36780 40588
rect 33600 40468 33652 40477
rect 33876 40400 33928 40452
rect 35716 40468 35768 40520
rect 36636 40468 36688 40520
rect 37004 40511 37056 40520
rect 37004 40477 37013 40511
rect 37013 40477 37047 40511
rect 37047 40477 37056 40511
rect 38108 40511 38160 40520
rect 37004 40468 37056 40477
rect 38108 40477 38117 40511
rect 38117 40477 38151 40511
rect 38151 40477 38160 40511
rect 38108 40468 38160 40477
rect 38200 40511 38252 40520
rect 38200 40477 38209 40511
rect 38209 40477 38243 40511
rect 38243 40477 38252 40511
rect 42984 40579 43036 40588
rect 42984 40545 42993 40579
rect 42993 40545 43027 40579
rect 43027 40545 43036 40579
rect 42984 40536 43036 40545
rect 46296 40579 46348 40588
rect 38200 40468 38252 40477
rect 40224 40511 40276 40520
rect 40224 40477 40233 40511
rect 40233 40477 40267 40511
rect 40267 40477 40276 40511
rect 40224 40468 40276 40477
rect 42524 40468 42576 40520
rect 43812 40511 43864 40520
rect 43812 40477 43821 40511
rect 43821 40477 43855 40511
rect 43855 40477 43864 40511
rect 43812 40468 43864 40477
rect 46296 40545 46305 40579
rect 46305 40545 46339 40579
rect 46339 40545 46348 40579
rect 46296 40536 46348 40545
rect 37372 40443 37424 40452
rect 37372 40409 37381 40443
rect 37381 40409 37415 40443
rect 37415 40409 37424 40443
rect 37556 40443 37608 40452
rect 37372 40400 37424 40409
rect 37556 40409 37565 40443
rect 37565 40409 37599 40443
rect 37599 40409 37608 40443
rect 37556 40400 37608 40409
rect 40684 40400 40736 40452
rect 46940 40400 46992 40452
rect 48136 40443 48188 40452
rect 48136 40409 48145 40443
rect 48145 40409 48179 40443
rect 48179 40409 48188 40443
rect 48136 40400 48188 40409
rect 28172 40375 28224 40384
rect 28172 40341 28181 40375
rect 28181 40341 28215 40375
rect 28215 40341 28224 40375
rect 28172 40332 28224 40341
rect 30748 40332 30800 40384
rect 35348 40375 35400 40384
rect 35348 40341 35357 40375
rect 35357 40341 35391 40375
rect 35391 40341 35400 40375
rect 35348 40332 35400 40341
rect 36360 40375 36412 40384
rect 36360 40341 36369 40375
rect 36369 40341 36403 40375
rect 36403 40341 36412 40375
rect 36360 40332 36412 40341
rect 36544 40332 36596 40384
rect 37464 40332 37516 40384
rect 41236 40332 41288 40384
rect 42524 40375 42576 40384
rect 42524 40341 42533 40375
rect 42533 40341 42567 40375
rect 42567 40341 42576 40375
rect 42524 40332 42576 40341
rect 42984 40332 43036 40384
rect 44180 40375 44232 40384
rect 44180 40341 44189 40375
rect 44189 40341 44223 40375
rect 44223 40341 44232 40375
rect 44180 40332 44232 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 23848 40128 23900 40180
rect 23480 40060 23532 40112
rect 24400 40060 24452 40112
rect 27988 40128 28040 40180
rect 35900 40128 35952 40180
rect 37556 40128 37608 40180
rect 44088 40128 44140 40180
rect 44732 40128 44784 40180
rect 27252 40060 27304 40112
rect 23664 39831 23716 39840
rect 23664 39797 23673 39831
rect 23673 39797 23707 39831
rect 23707 39797 23716 39831
rect 23664 39788 23716 39797
rect 24860 39788 24912 39840
rect 29552 40060 29604 40112
rect 29184 40035 29236 40044
rect 29184 40001 29193 40035
rect 29193 40001 29227 40035
rect 29227 40001 29236 40035
rect 29184 39992 29236 40001
rect 30196 40035 30248 40044
rect 30196 40001 30205 40035
rect 30205 40001 30239 40035
rect 30239 40001 30248 40035
rect 30196 39992 30248 40001
rect 31760 39992 31812 40044
rect 44180 40060 44232 40112
rect 45836 39992 45888 40044
rect 43996 39924 44048 39976
rect 31024 39856 31076 39908
rect 46940 40035 46992 40044
rect 46940 40001 46949 40035
rect 46949 40001 46983 40035
rect 46983 40001 46992 40035
rect 46940 39992 46992 40001
rect 27896 39788 27948 39840
rect 30012 39831 30064 39840
rect 30012 39797 30021 39831
rect 30021 39797 30055 39831
rect 30055 39797 30064 39831
rect 30012 39788 30064 39797
rect 47768 39831 47820 39840
rect 47768 39797 47777 39831
rect 47777 39797 47811 39831
rect 47811 39797 47820 39831
rect 47768 39788 47820 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 26608 39627 26660 39636
rect 26608 39593 26617 39627
rect 26617 39593 26651 39627
rect 26651 39593 26660 39627
rect 26608 39584 26660 39593
rect 27068 39584 27120 39636
rect 32588 39627 32640 39636
rect 32588 39593 32597 39627
rect 32597 39593 32631 39627
rect 32631 39593 32640 39627
rect 32588 39584 32640 39593
rect 38568 39584 38620 39636
rect 45100 39584 45152 39636
rect 27988 39516 28040 39568
rect 27068 39380 27120 39432
rect 27896 39423 27948 39432
rect 27896 39389 27905 39423
rect 27905 39389 27939 39423
rect 27939 39389 27948 39423
rect 27896 39380 27948 39389
rect 30196 39380 30248 39432
rect 30748 39423 30800 39432
rect 30748 39389 30757 39423
rect 30757 39389 30791 39423
rect 30791 39389 30800 39423
rect 30748 39380 30800 39389
rect 30840 39423 30892 39432
rect 30840 39389 30849 39423
rect 30849 39389 30883 39423
rect 30883 39389 30892 39423
rect 30840 39380 30892 39389
rect 31760 39380 31812 39432
rect 36636 39516 36688 39568
rect 34796 39380 34848 39432
rect 35900 39448 35952 39500
rect 39120 39448 39172 39500
rect 42800 39448 42852 39500
rect 47768 39448 47820 39500
rect 35348 39380 35400 39432
rect 35440 39423 35492 39432
rect 35440 39389 35449 39423
rect 35449 39389 35483 39423
rect 35483 39389 35492 39423
rect 35440 39380 35492 39389
rect 42524 39380 42576 39432
rect 42984 39423 43036 39432
rect 42984 39389 42993 39423
rect 42993 39389 43027 39423
rect 43027 39389 43036 39423
rect 42984 39380 43036 39389
rect 23664 39312 23716 39364
rect 24860 39312 24912 39364
rect 27712 39312 27764 39364
rect 39304 39312 39356 39364
rect 40408 39312 40460 39364
rect 25688 39244 25740 39296
rect 27804 39287 27856 39296
rect 27804 39253 27813 39287
rect 27813 39253 27847 39287
rect 27847 39253 27856 39287
rect 27804 39244 27856 39253
rect 28540 39244 28592 39296
rect 31484 39287 31536 39296
rect 31484 39253 31493 39287
rect 31493 39253 31527 39287
rect 31527 39253 31536 39287
rect 31484 39244 31536 39253
rect 34796 39287 34848 39296
rect 34796 39253 34805 39287
rect 34805 39253 34839 39287
rect 34839 39253 34848 39287
rect 34796 39244 34848 39253
rect 42340 39312 42392 39364
rect 47676 39312 47728 39364
rect 48136 39355 48188 39364
rect 48136 39321 48145 39355
rect 48145 39321 48179 39355
rect 48179 39321 48188 39355
rect 48136 39312 48188 39321
rect 42708 39244 42760 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 24584 39040 24636 39092
rect 31024 39040 31076 39092
rect 35440 39040 35492 39092
rect 41052 39083 41104 39092
rect 30840 38972 30892 39024
rect 30012 38947 30064 38956
rect 30012 38913 30021 38947
rect 30021 38913 30055 38947
rect 30055 38913 30064 38947
rect 31852 38972 31904 39024
rect 30012 38904 30064 38913
rect 40408 38972 40460 39024
rect 39120 38947 39172 38956
rect 30196 38836 30248 38888
rect 30932 38836 30984 38888
rect 31760 38836 31812 38888
rect 32220 38836 32272 38888
rect 33692 38879 33744 38888
rect 33692 38845 33701 38879
rect 33701 38845 33735 38879
rect 33735 38845 33744 38879
rect 33692 38836 33744 38845
rect 35348 38836 35400 38888
rect 37096 38836 37148 38888
rect 39120 38913 39129 38947
rect 39129 38913 39163 38947
rect 39163 38913 39172 38947
rect 39120 38904 39172 38913
rect 39304 38947 39356 38956
rect 39304 38913 39313 38947
rect 39313 38913 39347 38947
rect 39347 38913 39356 38947
rect 39304 38904 39356 38913
rect 37832 38836 37884 38888
rect 38200 38811 38252 38820
rect 38200 38777 38209 38811
rect 38209 38777 38243 38811
rect 38243 38777 38252 38811
rect 38200 38768 38252 38777
rect 41052 39049 41061 39083
rect 41061 39049 41095 39083
rect 41095 39049 41104 39083
rect 41052 39040 41104 39049
rect 41880 39040 41932 39092
rect 47676 39083 47728 39092
rect 47676 39049 47685 39083
rect 47685 39049 47719 39083
rect 47719 39049 47728 39083
rect 47676 39040 47728 39049
rect 41420 38972 41472 39024
rect 42708 38947 42760 38956
rect 42708 38913 42742 38947
rect 42742 38913 42760 38947
rect 42708 38904 42760 38913
rect 43996 38904 44048 38956
rect 40592 38768 40644 38820
rect 40776 38811 40828 38820
rect 40776 38777 40785 38811
rect 40785 38777 40819 38811
rect 40819 38777 40828 38811
rect 40776 38768 40828 38777
rect 41788 38768 41840 38820
rect 29828 38700 29880 38752
rect 32864 38700 32916 38752
rect 35624 38700 35676 38752
rect 38936 38743 38988 38752
rect 38936 38709 38945 38743
rect 38945 38709 38979 38743
rect 38979 38709 38988 38743
rect 38936 38700 38988 38709
rect 40132 38700 40184 38752
rect 41420 38700 41472 38752
rect 42156 38700 42208 38752
rect 46756 38904 46808 38956
rect 47584 38947 47636 38956
rect 47584 38913 47593 38947
rect 47593 38913 47627 38947
rect 47627 38913 47636 38947
rect 47584 38904 47636 38913
rect 45560 38700 45612 38752
rect 46572 38743 46624 38752
rect 46572 38709 46581 38743
rect 46581 38709 46615 38743
rect 46615 38709 46624 38743
rect 46572 38700 46624 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 26056 38496 26108 38548
rect 40960 38496 41012 38548
rect 41052 38496 41104 38548
rect 41604 38496 41656 38548
rect 42064 38539 42116 38548
rect 42064 38505 42073 38539
rect 42073 38505 42107 38539
rect 42107 38505 42116 38539
rect 42340 38539 42392 38548
rect 42064 38496 42116 38505
rect 42340 38505 42349 38539
rect 42349 38505 42383 38539
rect 42383 38505 42392 38539
rect 42340 38496 42392 38505
rect 46756 38539 46808 38548
rect 46756 38505 46765 38539
rect 46765 38505 46799 38539
rect 46799 38505 46808 38539
rect 46756 38496 46808 38505
rect 32220 38471 32272 38480
rect 32220 38437 32229 38471
rect 32229 38437 32263 38471
rect 32263 38437 32272 38471
rect 32220 38428 32272 38437
rect 29552 38360 29604 38412
rect 33692 38360 33744 38412
rect 42064 38403 42116 38412
rect 42064 38369 42073 38403
rect 42073 38369 42107 38403
rect 42107 38369 42116 38403
rect 45928 38403 45980 38412
rect 42064 38360 42116 38369
rect 45928 38369 45937 38403
rect 45937 38369 45971 38403
rect 45971 38369 45980 38403
rect 45928 38360 45980 38369
rect 46572 38360 46624 38412
rect 25780 38335 25832 38344
rect 25780 38301 25789 38335
rect 25789 38301 25823 38335
rect 25823 38301 25832 38335
rect 25780 38292 25832 38301
rect 28172 38292 28224 38344
rect 30748 38292 30800 38344
rect 32128 38292 32180 38344
rect 32864 38335 32916 38344
rect 32864 38301 32873 38335
rect 32873 38301 32907 38335
rect 32907 38301 32916 38335
rect 32864 38292 32916 38301
rect 34796 38292 34848 38344
rect 37188 38335 37240 38344
rect 37188 38301 37197 38335
rect 37197 38301 37231 38335
rect 37231 38301 37240 38335
rect 37188 38292 37240 38301
rect 38200 38292 38252 38344
rect 29736 38224 29788 38276
rect 25596 38199 25648 38208
rect 25596 38165 25605 38199
rect 25605 38165 25639 38199
rect 25639 38165 25648 38199
rect 25596 38156 25648 38165
rect 28908 38199 28960 38208
rect 28908 38165 28917 38199
rect 28917 38165 28951 38199
rect 28951 38165 28960 38199
rect 28908 38156 28960 38165
rect 30104 38199 30156 38208
rect 30104 38165 30113 38199
rect 30113 38165 30147 38199
rect 30147 38165 30156 38199
rect 30104 38156 30156 38165
rect 30196 38199 30248 38208
rect 30196 38165 30205 38199
rect 30205 38165 30239 38199
rect 30239 38165 30248 38199
rect 31484 38224 31536 38276
rect 30196 38156 30248 38165
rect 31300 38156 31352 38208
rect 32220 38156 32272 38208
rect 32680 38199 32732 38208
rect 32680 38165 32689 38199
rect 32689 38165 32723 38199
rect 32723 38165 32732 38199
rect 32680 38156 32732 38165
rect 35348 38156 35400 38208
rect 36452 38156 36504 38208
rect 40776 38292 40828 38344
rect 42800 38292 42852 38344
rect 43904 38292 43956 38344
rect 45100 38335 45152 38344
rect 45100 38301 45109 38335
rect 45109 38301 45143 38335
rect 45143 38301 45152 38335
rect 45100 38292 45152 38301
rect 47400 38335 47452 38344
rect 41512 38224 41564 38276
rect 41880 38267 41932 38276
rect 41880 38233 41889 38267
rect 41889 38233 41923 38267
rect 41923 38233 41932 38267
rect 41880 38224 41932 38233
rect 43812 38224 43864 38276
rect 44088 38224 44140 38276
rect 47400 38301 47409 38335
rect 47409 38301 47443 38335
rect 47443 38301 47452 38335
rect 47400 38292 47452 38301
rect 40224 38156 40276 38208
rect 40500 38156 40552 38208
rect 41604 38156 41656 38208
rect 42064 38156 42116 38208
rect 45100 38156 45152 38208
rect 46296 38199 46348 38208
rect 46296 38165 46305 38199
rect 46305 38165 46339 38199
rect 46339 38165 46348 38199
rect 46296 38156 46348 38165
rect 47492 38199 47544 38208
rect 47492 38165 47501 38199
rect 47501 38165 47535 38199
rect 47535 38165 47544 38199
rect 47492 38156 47544 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 30104 37952 30156 38004
rect 35624 37995 35676 38004
rect 24860 37748 24912 37800
rect 27620 37884 27672 37936
rect 25596 37816 25648 37868
rect 30196 37884 30248 37936
rect 29460 37859 29512 37868
rect 29460 37825 29494 37859
rect 29494 37825 29512 37859
rect 29460 37816 29512 37825
rect 29736 37816 29788 37868
rect 35624 37961 35633 37995
rect 35633 37961 35667 37995
rect 35667 37961 35676 37995
rect 35624 37952 35676 37961
rect 32680 37884 32732 37936
rect 37096 37952 37148 38004
rect 40776 37952 40828 38004
rect 41788 37995 41840 38004
rect 41788 37961 41797 37995
rect 41797 37961 41831 37995
rect 41831 37961 41840 37995
rect 41788 37952 41840 37961
rect 43812 37952 43864 38004
rect 31300 37859 31352 37868
rect 31300 37825 31309 37859
rect 31309 37825 31343 37859
rect 31343 37825 31352 37859
rect 35716 37859 35768 37868
rect 31300 37816 31352 37825
rect 35716 37825 35725 37859
rect 35725 37825 35759 37859
rect 35759 37825 35768 37859
rect 36452 37859 36504 37868
rect 35716 37816 35768 37825
rect 36452 37825 36461 37859
rect 36461 37825 36495 37859
rect 36495 37825 36504 37859
rect 36452 37816 36504 37825
rect 32128 37791 32180 37800
rect 26792 37612 26844 37664
rect 30748 37612 30800 37664
rect 32128 37757 32137 37791
rect 32137 37757 32171 37791
rect 32171 37757 32180 37791
rect 32128 37748 32180 37757
rect 35348 37791 35400 37800
rect 35348 37757 35357 37791
rect 35357 37757 35391 37791
rect 35391 37757 35400 37791
rect 35348 37748 35400 37757
rect 35624 37748 35676 37800
rect 37188 37816 37240 37868
rect 35992 37655 36044 37664
rect 35992 37621 36001 37655
rect 36001 37621 36035 37655
rect 36035 37621 36044 37655
rect 35992 37612 36044 37621
rect 36268 37612 36320 37664
rect 38936 37816 38988 37868
rect 40132 37816 40184 37868
rect 41420 37859 41472 37868
rect 41420 37825 41429 37859
rect 41429 37825 41463 37859
rect 41463 37825 41472 37859
rect 41420 37816 41472 37825
rect 40960 37748 41012 37800
rect 44272 37816 44324 37868
rect 45560 37816 45612 37868
rect 46296 37816 46348 37868
rect 40500 37612 40552 37664
rect 46940 37612 46992 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 25780 37408 25832 37460
rect 29460 37408 29512 37460
rect 41512 37451 41564 37460
rect 41512 37417 41521 37451
rect 41521 37417 41555 37451
rect 41555 37417 41564 37451
rect 41512 37408 41564 37417
rect 26792 37315 26844 37324
rect 26792 37281 26801 37315
rect 26801 37281 26835 37315
rect 26835 37281 26844 37315
rect 26792 37272 26844 37281
rect 27068 37272 27120 37324
rect 29552 37340 29604 37392
rect 29000 37315 29052 37324
rect 24952 37247 25004 37256
rect 24952 37213 24961 37247
rect 24961 37213 24995 37247
rect 24995 37213 25004 37247
rect 24952 37204 25004 37213
rect 25780 37247 25832 37256
rect 25780 37213 25789 37247
rect 25789 37213 25823 37247
rect 25823 37213 25832 37247
rect 25780 37204 25832 37213
rect 26976 37247 27028 37256
rect 26976 37213 26985 37247
rect 26985 37213 27019 37247
rect 27019 37213 27028 37247
rect 26976 37204 27028 37213
rect 28540 37247 28592 37256
rect 28540 37213 28549 37247
rect 28549 37213 28583 37247
rect 28583 37213 28592 37247
rect 28540 37204 28592 37213
rect 29000 37281 29009 37315
rect 29009 37281 29043 37315
rect 29043 37281 29052 37315
rect 29000 37272 29052 37281
rect 35624 37340 35676 37392
rect 36452 37340 36504 37392
rect 35348 37272 35400 37324
rect 41880 37340 41932 37392
rect 42248 37340 42300 37392
rect 44088 37340 44140 37392
rect 40776 37272 40828 37324
rect 28908 37204 28960 37256
rect 29828 37247 29880 37256
rect 29828 37213 29837 37247
rect 29837 37213 29871 37247
rect 29871 37213 29880 37247
rect 29828 37204 29880 37213
rect 35716 37204 35768 37256
rect 36452 37247 36504 37256
rect 36452 37213 36461 37247
rect 36461 37213 36495 37247
rect 36495 37213 36504 37247
rect 36452 37204 36504 37213
rect 37096 37204 37148 37256
rect 40960 37204 41012 37256
rect 28724 37179 28776 37188
rect 28724 37145 28733 37179
rect 28733 37145 28767 37179
rect 28767 37145 28776 37179
rect 28724 37136 28776 37145
rect 30932 37136 30984 37188
rect 31852 37136 31904 37188
rect 43996 37247 44048 37256
rect 43996 37213 44005 37247
rect 44005 37213 44039 37247
rect 44039 37213 44048 37247
rect 43996 37204 44048 37213
rect 44272 37247 44324 37256
rect 43812 37136 43864 37188
rect 44272 37213 44281 37247
rect 44281 37213 44315 37247
rect 44315 37213 44324 37247
rect 44272 37204 44324 37213
rect 46296 37247 46348 37256
rect 46296 37213 46305 37247
rect 46305 37213 46339 37247
rect 46339 37213 46348 37247
rect 46296 37204 46348 37213
rect 47492 37136 47544 37188
rect 48136 37179 48188 37188
rect 48136 37145 48145 37179
rect 48145 37145 48179 37179
rect 48179 37145 48188 37179
rect 48136 37136 48188 37145
rect 24676 37068 24728 37120
rect 27252 37068 27304 37120
rect 28356 37111 28408 37120
rect 28356 37077 28365 37111
rect 28365 37077 28399 37111
rect 28399 37077 28408 37111
rect 28356 37068 28408 37077
rect 35440 37068 35492 37120
rect 36360 37068 36412 37120
rect 36912 37111 36964 37120
rect 36912 37077 36921 37111
rect 36921 37077 36955 37111
rect 36955 37077 36964 37111
rect 36912 37068 36964 37077
rect 41420 37068 41472 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 36912 36864 36964 36916
rect 24308 36771 24360 36780
rect 24308 36737 24342 36771
rect 24342 36737 24360 36771
rect 27620 36796 27672 36848
rect 27896 36796 27948 36848
rect 28356 36796 28408 36848
rect 44732 36839 44784 36848
rect 24308 36728 24360 36737
rect 27252 36771 27304 36780
rect 27252 36737 27286 36771
rect 27286 36737 27304 36771
rect 27252 36728 27304 36737
rect 33140 36771 33192 36780
rect 33140 36737 33174 36771
rect 33174 36737 33192 36771
rect 33140 36728 33192 36737
rect 31760 36660 31812 36712
rect 32128 36660 32180 36712
rect 44732 36805 44741 36839
rect 44741 36805 44775 36839
rect 44775 36805 44784 36839
rect 44732 36796 44784 36805
rect 46204 36796 46256 36848
rect 46296 36796 46348 36848
rect 35992 36771 36044 36780
rect 24400 36524 24452 36576
rect 24768 36524 24820 36576
rect 25412 36567 25464 36576
rect 25412 36533 25421 36567
rect 25421 36533 25455 36567
rect 25455 36533 25464 36567
rect 25412 36524 25464 36533
rect 27160 36524 27212 36576
rect 30196 36567 30248 36576
rect 30196 36533 30205 36567
rect 30205 36533 30239 36567
rect 30239 36533 30248 36567
rect 30196 36524 30248 36533
rect 34244 36567 34296 36576
rect 34244 36533 34253 36567
rect 34253 36533 34287 36567
rect 34287 36533 34296 36567
rect 34244 36524 34296 36533
rect 34520 36524 34572 36576
rect 35992 36737 36001 36771
rect 36001 36737 36035 36771
rect 36035 36737 36044 36771
rect 35992 36728 36044 36737
rect 36268 36771 36320 36780
rect 36268 36737 36277 36771
rect 36277 36737 36311 36771
rect 36311 36737 36320 36771
rect 36268 36728 36320 36737
rect 39856 36728 39908 36780
rect 41420 36771 41472 36780
rect 41420 36737 41429 36771
rect 41429 36737 41463 36771
rect 41463 36737 41472 36771
rect 47032 36771 47084 36780
rect 41420 36728 41472 36737
rect 47032 36737 47041 36771
rect 47041 36737 47075 36771
rect 47075 36737 47084 36771
rect 47032 36728 47084 36737
rect 35624 36592 35676 36644
rect 35348 36524 35400 36576
rect 36268 36592 36320 36644
rect 40408 36592 40460 36644
rect 43996 36592 44048 36644
rect 44180 36592 44232 36644
rect 35808 36567 35860 36576
rect 35808 36533 35817 36567
rect 35817 36533 35851 36567
rect 35851 36533 35860 36567
rect 40500 36567 40552 36576
rect 35808 36524 35860 36533
rect 40500 36533 40509 36567
rect 40509 36533 40543 36567
rect 40543 36533 40552 36567
rect 40500 36524 40552 36533
rect 41236 36567 41288 36576
rect 41236 36533 41245 36567
rect 41245 36533 41279 36567
rect 41279 36533 41288 36567
rect 41236 36524 41288 36533
rect 45192 36524 45244 36576
rect 45836 36524 45888 36576
rect 46664 36524 46716 36576
rect 46848 36567 46900 36576
rect 46848 36533 46857 36567
rect 46857 36533 46891 36567
rect 46891 36533 46900 36567
rect 46848 36524 46900 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 25780 36363 25832 36372
rect 25780 36329 25789 36363
rect 25789 36329 25823 36363
rect 25823 36329 25832 36363
rect 25780 36320 25832 36329
rect 26884 36320 26936 36372
rect 42248 36363 42300 36372
rect 27252 36252 27304 36304
rect 40408 36295 40460 36304
rect 40408 36261 40417 36295
rect 40417 36261 40451 36295
rect 40451 36261 40460 36295
rect 40408 36252 40460 36261
rect 42248 36329 42257 36363
rect 42257 36329 42291 36363
rect 42291 36329 42300 36363
rect 42248 36320 42300 36329
rect 45836 36320 45888 36372
rect 46204 36320 46256 36372
rect 46940 36320 46992 36372
rect 29184 36184 29236 36236
rect 30196 36184 30248 36236
rect 34244 36184 34296 36236
rect 36452 36227 36504 36236
rect 36452 36193 36461 36227
rect 36461 36193 36495 36227
rect 36495 36193 36504 36227
rect 36452 36184 36504 36193
rect 45560 36184 45612 36236
rect 46756 36227 46808 36236
rect 46756 36193 46765 36227
rect 46765 36193 46799 36227
rect 46799 36193 46808 36227
rect 46756 36184 46808 36193
rect 19984 36116 20036 36168
rect 24400 36159 24452 36168
rect 24400 36125 24409 36159
rect 24409 36125 24443 36159
rect 24443 36125 24452 36159
rect 24400 36116 24452 36125
rect 24676 36159 24728 36168
rect 24676 36125 24710 36159
rect 24710 36125 24728 36159
rect 24676 36116 24728 36125
rect 26792 36116 26844 36168
rect 27160 36116 27212 36168
rect 27344 36116 27396 36168
rect 30932 36116 30984 36168
rect 34980 36159 35032 36168
rect 34980 36125 34989 36159
rect 34989 36125 35023 36159
rect 35023 36125 35032 36159
rect 34980 36116 35032 36125
rect 35440 36116 35492 36168
rect 36268 36159 36320 36168
rect 36268 36125 36277 36159
rect 36277 36125 36311 36159
rect 36311 36125 36320 36159
rect 36268 36116 36320 36125
rect 26700 36048 26752 36100
rect 20444 35980 20496 36032
rect 26884 35980 26936 36032
rect 35624 36048 35676 36100
rect 36912 36116 36964 36168
rect 42800 36116 42852 36168
rect 45928 36159 45980 36168
rect 45928 36125 45937 36159
rect 45937 36125 45971 36159
rect 45971 36125 45980 36159
rect 45928 36116 45980 36125
rect 46848 36116 46900 36168
rect 40960 36048 41012 36100
rect 41236 36048 41288 36100
rect 42984 36091 43036 36100
rect 42984 36057 43018 36091
rect 43018 36057 43036 36091
rect 42984 36048 43036 36057
rect 46572 36048 46624 36100
rect 27804 35980 27856 36032
rect 29552 35980 29604 36032
rect 35992 36023 36044 36032
rect 35992 35989 36001 36023
rect 36001 35989 36035 36023
rect 36035 35989 36044 36023
rect 35992 35980 36044 35989
rect 44088 36023 44140 36032
rect 44088 35989 44097 36023
rect 44097 35989 44131 36023
rect 44131 35989 44140 36023
rect 44088 35980 44140 35989
rect 46388 35980 46440 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 24308 35776 24360 35828
rect 24952 35776 25004 35828
rect 37004 35776 37056 35828
rect 40684 35819 40736 35828
rect 40684 35785 40693 35819
rect 40693 35785 40727 35819
rect 40727 35785 40736 35819
rect 40684 35776 40736 35785
rect 42984 35776 43036 35828
rect 44088 35776 44140 35828
rect 26056 35708 26108 35760
rect 27068 35708 27120 35760
rect 24952 35640 25004 35692
rect 25044 35683 25096 35692
rect 25044 35649 25053 35683
rect 25053 35649 25087 35683
rect 25087 35649 25096 35683
rect 25044 35640 25096 35649
rect 25872 35640 25924 35692
rect 27252 35683 27304 35692
rect 27252 35649 27261 35683
rect 27261 35649 27295 35683
rect 27295 35649 27304 35683
rect 27252 35640 27304 35649
rect 29552 35683 29604 35692
rect 29552 35649 29561 35683
rect 29561 35649 29595 35683
rect 29595 35649 29604 35683
rect 29552 35640 29604 35649
rect 32312 35683 32364 35692
rect 32312 35649 32321 35683
rect 32321 35649 32355 35683
rect 32355 35649 32364 35683
rect 32312 35640 32364 35649
rect 33508 35640 33560 35692
rect 34980 35640 35032 35692
rect 35256 35683 35308 35692
rect 35256 35649 35265 35683
rect 35265 35649 35299 35683
rect 35299 35649 35308 35683
rect 35256 35640 35308 35649
rect 36452 35708 36504 35760
rect 43996 35751 44048 35760
rect 43996 35717 44005 35751
rect 44005 35717 44039 35751
rect 44039 35717 44048 35751
rect 43996 35708 44048 35717
rect 44364 35708 44416 35760
rect 35440 35683 35492 35692
rect 35440 35649 35449 35683
rect 35449 35649 35483 35683
rect 35483 35649 35492 35683
rect 35440 35640 35492 35649
rect 35624 35683 35676 35692
rect 35624 35649 35633 35683
rect 35633 35649 35667 35683
rect 35667 35649 35676 35683
rect 38936 35683 38988 35692
rect 35624 35640 35676 35649
rect 38936 35649 38945 35683
rect 38945 35649 38979 35683
rect 38979 35649 38988 35683
rect 38936 35640 38988 35649
rect 39948 35683 40000 35692
rect 39948 35649 39957 35683
rect 39957 35649 39991 35683
rect 39991 35649 40000 35683
rect 40868 35683 40920 35692
rect 39948 35640 40000 35649
rect 40868 35649 40877 35683
rect 40877 35649 40911 35683
rect 40911 35649 40920 35683
rect 40868 35640 40920 35649
rect 42984 35683 43036 35692
rect 42984 35649 42993 35683
rect 42993 35649 43027 35683
rect 43027 35649 43036 35683
rect 42984 35640 43036 35649
rect 44640 35640 44692 35692
rect 47032 35776 47084 35828
rect 45744 35683 45796 35692
rect 45744 35649 45753 35683
rect 45753 35649 45787 35683
rect 45787 35649 45796 35683
rect 45744 35640 45796 35649
rect 46388 35683 46440 35692
rect 46388 35649 46397 35683
rect 46397 35649 46431 35683
rect 46431 35649 46440 35683
rect 46388 35640 46440 35649
rect 46940 35640 46992 35692
rect 47768 35683 47820 35692
rect 47768 35649 47777 35683
rect 47777 35649 47811 35683
rect 47811 35649 47820 35683
rect 47768 35640 47820 35649
rect 25412 35572 25464 35624
rect 25504 35572 25556 35624
rect 27160 35615 27212 35624
rect 27160 35581 27169 35615
rect 27169 35581 27203 35615
rect 27203 35581 27212 35615
rect 27160 35572 27212 35581
rect 33232 35572 33284 35624
rect 38568 35572 38620 35624
rect 43720 35615 43772 35624
rect 43720 35581 43729 35615
rect 43729 35581 43763 35615
rect 43763 35581 43772 35615
rect 43720 35572 43772 35581
rect 44180 35572 44232 35624
rect 26792 35504 26844 35556
rect 25688 35436 25740 35488
rect 25964 35479 26016 35488
rect 25964 35445 25973 35479
rect 25973 35445 26007 35479
rect 26007 35445 26016 35479
rect 25964 35436 26016 35445
rect 26148 35479 26200 35488
rect 26148 35445 26157 35479
rect 26157 35445 26191 35479
rect 26191 35445 26200 35479
rect 26148 35436 26200 35445
rect 28724 35504 28776 35556
rect 32128 35504 32180 35556
rect 40408 35504 40460 35556
rect 45192 35572 45244 35624
rect 46572 35615 46624 35624
rect 46572 35581 46581 35615
rect 46581 35581 46615 35615
rect 46615 35581 46624 35615
rect 46572 35572 46624 35581
rect 27068 35436 27120 35488
rect 29000 35436 29052 35488
rect 29368 35479 29420 35488
rect 29368 35445 29377 35479
rect 29377 35445 29411 35479
rect 29411 35445 29420 35479
rect 29368 35436 29420 35445
rect 32220 35436 32272 35488
rect 34704 35436 34756 35488
rect 37372 35436 37424 35488
rect 40132 35436 40184 35488
rect 43444 35479 43496 35488
rect 43444 35445 43453 35479
rect 43453 35445 43487 35479
rect 43487 35445 43496 35479
rect 43444 35436 43496 35445
rect 44732 35436 44784 35488
rect 46020 35436 46072 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 24952 35232 25004 35284
rect 33416 35232 33468 35284
rect 38660 35232 38712 35284
rect 26056 35096 26108 35148
rect 42984 35232 43036 35284
rect 46572 35232 46624 35284
rect 2044 35028 2096 35080
rect 25044 35071 25096 35080
rect 25044 35037 25053 35071
rect 25053 35037 25087 35071
rect 25087 35037 25096 35071
rect 25044 35028 25096 35037
rect 25504 35028 25556 35080
rect 27804 35071 27856 35080
rect 27804 35037 27813 35071
rect 27813 35037 27847 35071
rect 27847 35037 27856 35071
rect 27804 35028 27856 35037
rect 29000 35028 29052 35080
rect 31760 35028 31812 35080
rect 34704 35071 34756 35080
rect 34704 35037 34713 35071
rect 34713 35037 34747 35071
rect 34747 35037 34756 35071
rect 34704 35028 34756 35037
rect 34888 35071 34940 35080
rect 34888 35037 34897 35071
rect 34897 35037 34931 35071
rect 34931 35037 34940 35071
rect 34888 35028 34940 35037
rect 36176 35071 36228 35080
rect 36176 35037 36185 35071
rect 36185 35037 36219 35071
rect 36219 35037 36228 35071
rect 36176 35028 36228 35037
rect 24860 34960 24912 35012
rect 25872 35003 25924 35012
rect 25872 34969 25881 35003
rect 25881 34969 25915 35003
rect 25915 34969 25924 35003
rect 25872 34960 25924 34969
rect 25964 34892 26016 34944
rect 27528 34935 27580 34944
rect 27528 34901 27537 34935
rect 27537 34901 27571 34935
rect 27571 34901 27580 34935
rect 27528 34892 27580 34901
rect 27988 35003 28040 35012
rect 27988 34969 28023 35003
rect 28023 34969 28040 35003
rect 27988 34960 28040 34969
rect 32864 34960 32916 35012
rect 35900 35003 35952 35012
rect 35900 34969 35909 35003
rect 35909 34969 35943 35003
rect 35943 34969 35952 35003
rect 35900 34960 35952 34969
rect 39120 35096 39172 35148
rect 38936 35071 38988 35080
rect 38936 35037 38945 35071
rect 38945 35037 38979 35071
rect 38979 35037 38988 35071
rect 38936 35028 38988 35037
rect 43720 35096 43772 35148
rect 45744 35096 45796 35148
rect 46756 35139 46808 35148
rect 46756 35105 46765 35139
rect 46765 35105 46799 35139
rect 46799 35105 46808 35139
rect 46756 35096 46808 35105
rect 40500 35028 40552 35080
rect 44180 35028 44232 35080
rect 44732 35028 44784 35080
rect 40132 35003 40184 35012
rect 40132 34969 40166 35003
rect 40166 34969 40184 35003
rect 40132 34960 40184 34969
rect 46848 35028 46900 35080
rect 28724 34892 28776 34944
rect 32312 34935 32364 34944
rect 32312 34901 32321 34935
rect 32321 34901 32355 34935
rect 32355 34901 32364 34935
rect 32312 34892 32364 34901
rect 32680 34892 32732 34944
rect 34980 34892 35032 34944
rect 35440 34892 35492 34944
rect 37004 34892 37056 34944
rect 37280 34892 37332 34944
rect 38936 34892 38988 34944
rect 40224 34892 40276 34944
rect 45192 34892 45244 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 25412 34688 25464 34740
rect 25872 34688 25924 34740
rect 26148 34688 26200 34740
rect 27988 34688 28040 34740
rect 32864 34731 32916 34740
rect 32864 34697 32873 34731
rect 32873 34697 32907 34731
rect 32907 34697 32916 34731
rect 32864 34688 32916 34697
rect 34888 34688 34940 34740
rect 35900 34688 35952 34740
rect 39948 34688 40000 34740
rect 45744 34688 45796 34740
rect 46848 34731 46900 34740
rect 46848 34697 46857 34731
rect 46857 34697 46891 34731
rect 46891 34697 46900 34731
rect 46848 34688 46900 34697
rect 27528 34620 27580 34672
rect 29368 34620 29420 34672
rect 2044 34595 2096 34604
rect 2044 34561 2053 34595
rect 2053 34561 2087 34595
rect 2087 34561 2096 34595
rect 2044 34552 2096 34561
rect 24400 34595 24452 34604
rect 24400 34561 24409 34595
rect 24409 34561 24443 34595
rect 24443 34561 24452 34595
rect 24400 34552 24452 34561
rect 24492 34552 24544 34604
rect 27068 34595 27120 34604
rect 27068 34561 27077 34595
rect 27077 34561 27111 34595
rect 27111 34561 27120 34595
rect 27068 34552 27120 34561
rect 27896 34595 27948 34604
rect 27896 34561 27905 34595
rect 27905 34561 27939 34595
rect 27939 34561 27948 34595
rect 27896 34552 27948 34561
rect 32128 34595 32180 34604
rect 32128 34561 32137 34595
rect 32137 34561 32171 34595
rect 32171 34561 32180 34595
rect 32128 34552 32180 34561
rect 32312 34595 32364 34604
rect 32312 34561 32321 34595
rect 32321 34561 32355 34595
rect 32355 34561 32364 34595
rect 32312 34552 32364 34561
rect 32680 34595 32732 34604
rect 32680 34561 32689 34595
rect 32689 34561 32723 34595
rect 32723 34561 32732 34595
rect 32680 34552 32732 34561
rect 33416 34595 33468 34604
rect 33416 34561 33425 34595
rect 33425 34561 33459 34595
rect 33459 34561 33468 34595
rect 33416 34552 33468 34561
rect 33508 34552 33560 34604
rect 34612 34620 34664 34672
rect 43812 34620 43864 34672
rect 34428 34595 34480 34604
rect 34428 34561 34437 34595
rect 34437 34561 34471 34595
rect 34471 34561 34480 34595
rect 34428 34552 34480 34561
rect 34520 34595 34572 34604
rect 34520 34561 34529 34595
rect 34529 34561 34563 34595
rect 34563 34561 34572 34595
rect 34520 34552 34572 34561
rect 34704 34552 34756 34604
rect 34980 34595 35032 34604
rect 34980 34561 34989 34595
rect 34989 34561 35023 34595
rect 35023 34561 35032 34595
rect 34980 34552 35032 34561
rect 35348 34552 35400 34604
rect 35992 34552 36044 34604
rect 37004 34552 37056 34604
rect 37280 34595 37332 34604
rect 37280 34561 37289 34595
rect 37289 34561 37323 34595
rect 37323 34561 37332 34595
rect 37280 34552 37332 34561
rect 37372 34595 37424 34604
rect 37372 34561 37381 34595
rect 37381 34561 37415 34595
rect 37415 34561 37424 34595
rect 39028 34595 39080 34604
rect 37372 34552 37424 34561
rect 39028 34561 39037 34595
rect 39037 34561 39071 34595
rect 39071 34561 39080 34595
rect 39028 34552 39080 34561
rect 41144 34595 41196 34604
rect 41144 34561 41153 34595
rect 41153 34561 41187 34595
rect 41187 34561 41196 34595
rect 41144 34552 41196 34561
rect 42800 34552 42852 34604
rect 45008 34552 45060 34604
rect 46388 34552 46440 34604
rect 47768 34620 47820 34672
rect 2228 34527 2280 34536
rect 2228 34493 2237 34527
rect 2237 34493 2271 34527
rect 2271 34493 2280 34527
rect 2228 34484 2280 34493
rect 3608 34527 3660 34536
rect 3608 34493 3617 34527
rect 3617 34493 3651 34527
rect 3651 34493 3660 34527
rect 3608 34484 3660 34493
rect 29736 34527 29788 34536
rect 29736 34493 29745 34527
rect 29745 34493 29779 34527
rect 29779 34493 29788 34527
rect 29736 34484 29788 34493
rect 32128 34416 32180 34468
rect 33968 34484 34020 34536
rect 32956 34416 33008 34468
rect 38568 34484 38620 34536
rect 39120 34527 39172 34536
rect 39120 34493 39129 34527
rect 39129 34493 39163 34527
rect 39163 34493 39172 34527
rect 39120 34484 39172 34493
rect 41696 34484 41748 34536
rect 29276 34391 29328 34400
rect 29276 34357 29285 34391
rect 29285 34357 29319 34391
rect 29319 34357 29328 34391
rect 29276 34348 29328 34357
rect 31116 34391 31168 34400
rect 31116 34357 31125 34391
rect 31125 34357 31159 34391
rect 31159 34357 31168 34391
rect 31116 34348 31168 34357
rect 33324 34348 33376 34400
rect 34796 34348 34848 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 2228 34144 2280 34196
rect 24492 34144 24544 34196
rect 27620 34144 27672 34196
rect 27896 34144 27948 34196
rect 32312 34144 32364 34196
rect 32128 34119 32180 34128
rect 32128 34085 32137 34119
rect 32137 34085 32171 34119
rect 32171 34085 32180 34119
rect 32128 34076 32180 34085
rect 36176 34144 36228 34196
rect 40868 34144 40920 34196
rect 43812 34187 43864 34196
rect 43812 34153 43821 34187
rect 43821 34153 43855 34187
rect 43855 34153 43864 34187
rect 43812 34144 43864 34153
rect 45008 34187 45060 34196
rect 45008 34153 45017 34187
rect 45017 34153 45051 34187
rect 45051 34153 45060 34187
rect 45008 34144 45060 34153
rect 2412 33940 2464 33992
rect 18144 33940 18196 33992
rect 24860 33940 24912 33992
rect 30380 33940 30432 33992
rect 30656 33983 30708 33992
rect 30656 33949 30665 33983
rect 30665 33949 30699 33983
rect 30699 33949 30708 33983
rect 30656 33940 30708 33949
rect 31024 33940 31076 33992
rect 32128 33940 32180 33992
rect 32220 33940 32272 33992
rect 25964 33872 26016 33924
rect 28632 33872 28684 33924
rect 33416 34076 33468 34128
rect 37924 34008 37976 34060
rect 41696 34051 41748 34060
rect 41696 34017 41705 34051
rect 41705 34017 41739 34051
rect 41739 34017 41748 34051
rect 41696 34008 41748 34017
rect 46480 34008 46532 34060
rect 46756 34051 46808 34060
rect 46756 34017 46765 34051
rect 46765 34017 46799 34051
rect 46799 34017 46808 34051
rect 46756 34008 46808 34017
rect 33416 33940 33468 33992
rect 33968 33983 34020 33992
rect 33968 33949 33977 33983
rect 33977 33949 34011 33983
rect 34011 33949 34020 33983
rect 33968 33940 34020 33949
rect 34704 33983 34756 33992
rect 34704 33949 34713 33983
rect 34713 33949 34747 33983
rect 34747 33949 34756 33983
rect 34704 33940 34756 33949
rect 36360 33983 36412 33992
rect 36360 33949 36369 33983
rect 36369 33949 36403 33983
rect 36403 33949 36412 33983
rect 36360 33940 36412 33949
rect 40592 33940 40644 33992
rect 29000 33804 29052 33856
rect 34428 33872 34480 33924
rect 34520 33872 34572 33924
rect 34888 33915 34940 33924
rect 34888 33881 34897 33915
rect 34897 33881 34931 33915
rect 34931 33881 34940 33915
rect 34888 33872 34940 33881
rect 35348 33872 35400 33924
rect 41236 33940 41288 33992
rect 42892 33940 42944 33992
rect 43996 33983 44048 33992
rect 43996 33949 44005 33983
rect 44005 33949 44039 33983
rect 44039 33949 44048 33983
rect 43996 33940 44048 33949
rect 45192 33983 45244 33992
rect 45192 33949 45201 33983
rect 45201 33949 45235 33983
rect 45235 33949 45244 33983
rect 45192 33940 45244 33949
rect 43260 33872 43312 33924
rect 47676 33872 47728 33924
rect 32220 33804 32272 33856
rect 35072 33847 35124 33856
rect 35072 33813 35081 33847
rect 35081 33813 35115 33847
rect 35115 33813 35124 33847
rect 35072 33804 35124 33813
rect 48044 33804 48096 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 24400 33600 24452 33652
rect 25504 33643 25556 33652
rect 25504 33609 25513 33643
rect 25513 33609 25547 33643
rect 25547 33609 25556 33643
rect 25504 33600 25556 33609
rect 31208 33600 31260 33652
rect 30932 33575 30984 33584
rect 30932 33541 30941 33575
rect 30941 33541 30975 33575
rect 30975 33541 30984 33575
rect 30932 33532 30984 33541
rect 31024 33532 31076 33584
rect 26148 33507 26200 33516
rect 26148 33473 26157 33507
rect 26157 33473 26191 33507
rect 26191 33473 26200 33507
rect 26148 33464 26200 33473
rect 28632 33507 28684 33516
rect 28632 33473 28641 33507
rect 28641 33473 28675 33507
rect 28675 33473 28684 33507
rect 28632 33464 28684 33473
rect 31208 33464 31260 33516
rect 31668 33464 31720 33516
rect 33140 33532 33192 33584
rect 35072 33600 35124 33652
rect 41236 33643 41288 33652
rect 41236 33609 41245 33643
rect 41245 33609 41279 33643
rect 41279 33609 41288 33643
rect 41236 33600 41288 33609
rect 43260 33600 43312 33652
rect 42892 33532 42944 33584
rect 43444 33532 43496 33584
rect 33324 33464 33376 33516
rect 33508 33507 33560 33516
rect 33508 33473 33517 33507
rect 33517 33473 33551 33507
rect 33551 33473 33560 33507
rect 33508 33464 33560 33473
rect 29736 33396 29788 33448
rect 31760 33396 31812 33448
rect 32220 33396 32272 33448
rect 32588 33439 32640 33448
rect 32588 33405 32597 33439
rect 32597 33405 32631 33439
rect 32631 33405 32640 33439
rect 32588 33396 32640 33405
rect 33048 33396 33100 33448
rect 33876 33507 33928 33516
rect 33876 33473 33885 33507
rect 33885 33473 33919 33507
rect 33919 33473 33928 33507
rect 33876 33464 33928 33473
rect 34428 33464 34480 33516
rect 34796 33507 34848 33516
rect 34796 33473 34805 33507
rect 34805 33473 34839 33507
rect 34839 33473 34848 33507
rect 34796 33464 34848 33473
rect 41420 33507 41472 33516
rect 41420 33473 41429 33507
rect 41429 33473 41463 33507
rect 41463 33473 41472 33507
rect 42800 33507 42852 33516
rect 41420 33464 41472 33473
rect 42800 33473 42809 33507
rect 42809 33473 42843 33507
rect 42843 33473 42852 33507
rect 42800 33464 42852 33473
rect 44824 33507 44876 33516
rect 44824 33473 44833 33507
rect 44833 33473 44867 33507
rect 44867 33473 44876 33507
rect 44824 33464 44876 33473
rect 46848 33464 46900 33516
rect 38108 33328 38160 33380
rect 44732 33328 44784 33380
rect 32496 33260 32548 33312
rect 33232 33260 33284 33312
rect 35808 33260 35860 33312
rect 44640 33303 44692 33312
rect 44640 33269 44649 33303
rect 44649 33269 44683 33303
rect 44683 33269 44692 33303
rect 44640 33260 44692 33269
rect 46940 33260 46992 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 26148 33056 26200 33108
rect 30380 33099 30432 33108
rect 30380 33065 30389 33099
rect 30389 33065 30423 33099
rect 30423 33065 30432 33099
rect 30380 33056 30432 33065
rect 30656 33056 30708 33108
rect 31668 33099 31720 33108
rect 31668 33065 31677 33099
rect 31677 33065 31711 33099
rect 31711 33065 31720 33099
rect 31668 33056 31720 33065
rect 32588 33056 32640 33108
rect 33140 33056 33192 33108
rect 2136 32852 2188 32904
rect 24860 32920 24912 32972
rect 27620 32963 27672 32972
rect 25412 32895 25464 32904
rect 25412 32861 25421 32895
rect 25421 32861 25455 32895
rect 25455 32861 25464 32895
rect 25412 32852 25464 32861
rect 27620 32929 27629 32963
rect 27629 32929 27663 32963
rect 27663 32929 27672 32963
rect 27620 32920 27672 32929
rect 29276 32920 29328 32972
rect 29552 32920 29604 32972
rect 26056 32784 26108 32836
rect 25320 32716 25372 32768
rect 29000 32852 29052 32904
rect 32312 32988 32364 33040
rect 32496 32988 32548 33040
rect 34336 32988 34388 33040
rect 36360 33056 36412 33108
rect 38660 33056 38712 33108
rect 39764 33056 39816 33108
rect 40776 33099 40828 33108
rect 40776 33065 40785 33099
rect 40785 33065 40819 33099
rect 40819 33065 40828 33099
rect 40776 33056 40828 33065
rect 41420 33056 41472 33108
rect 42800 33056 42852 33108
rect 40132 32988 40184 33040
rect 41696 32988 41748 33040
rect 35900 32920 35952 32972
rect 44180 33056 44232 33108
rect 47676 33099 47728 33108
rect 31300 32895 31352 32904
rect 31300 32861 31309 32895
rect 31309 32861 31343 32895
rect 31343 32861 31352 32895
rect 31300 32852 31352 32861
rect 30380 32784 30432 32836
rect 31208 32784 31260 32836
rect 32404 32852 32456 32904
rect 33232 32895 33284 32904
rect 33232 32861 33241 32895
rect 33241 32861 33275 32895
rect 33275 32861 33284 32895
rect 33232 32852 33284 32861
rect 33416 32895 33468 32904
rect 33416 32861 33425 32895
rect 33425 32861 33459 32895
rect 33459 32861 33468 32895
rect 33416 32852 33468 32861
rect 33140 32784 33192 32836
rect 28816 32716 28868 32768
rect 32312 32716 32364 32768
rect 32496 32759 32548 32768
rect 32496 32725 32505 32759
rect 32505 32725 32539 32759
rect 32539 32725 32548 32759
rect 32496 32716 32548 32725
rect 32680 32716 32732 32768
rect 35808 32852 35860 32904
rect 37280 32852 37332 32904
rect 38016 32852 38068 32904
rect 43996 32895 44048 32904
rect 43996 32861 44005 32895
rect 44005 32861 44039 32895
rect 44039 32861 44048 32895
rect 43996 32852 44048 32861
rect 44640 32852 44692 32904
rect 47676 33065 47685 33099
rect 47685 33065 47719 33099
rect 47719 33065 47728 33099
rect 47676 33056 47728 33065
rect 35992 32784 36044 32836
rect 38568 32784 38620 32836
rect 40960 32784 41012 32836
rect 41604 32827 41656 32836
rect 41604 32793 41613 32827
rect 41613 32793 41647 32827
rect 41647 32793 41656 32827
rect 41604 32784 41656 32793
rect 40500 32716 40552 32768
rect 46112 32716 46164 32768
rect 47308 32784 47360 32836
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 2136 32419 2188 32428
rect 2136 32385 2145 32419
rect 2145 32385 2179 32419
rect 2179 32385 2188 32419
rect 2136 32376 2188 32385
rect 25320 32419 25372 32428
rect 25320 32385 25329 32419
rect 25329 32385 25363 32419
rect 25363 32385 25372 32419
rect 25320 32376 25372 32385
rect 29552 32512 29604 32564
rect 29736 32555 29788 32564
rect 29736 32521 29745 32555
rect 29745 32521 29779 32555
rect 29779 32521 29788 32555
rect 29736 32512 29788 32521
rect 32496 32555 32548 32564
rect 32496 32521 32505 32555
rect 32505 32521 32539 32555
rect 32539 32521 32548 32555
rect 32496 32512 32548 32521
rect 33140 32512 33192 32564
rect 34428 32512 34480 32564
rect 37096 32512 37148 32564
rect 37924 32555 37976 32564
rect 37924 32521 37933 32555
rect 37933 32521 37967 32555
rect 37967 32521 37976 32555
rect 37924 32512 37976 32521
rect 28816 32444 28868 32496
rect 29184 32376 29236 32428
rect 31668 32444 31720 32496
rect 33324 32444 33376 32496
rect 33416 32444 33468 32496
rect 34152 32444 34204 32496
rect 34336 32444 34388 32496
rect 30840 32419 30892 32428
rect 2504 32308 2556 32360
rect 2780 32351 2832 32360
rect 2780 32317 2789 32351
rect 2789 32317 2823 32351
rect 2823 32317 2832 32351
rect 2780 32308 2832 32317
rect 27620 32308 27672 32360
rect 28816 32351 28868 32360
rect 28816 32317 28825 32351
rect 28825 32317 28859 32351
rect 28859 32317 28868 32351
rect 28816 32308 28868 32317
rect 30840 32385 30849 32419
rect 30849 32385 30883 32419
rect 30883 32385 30892 32419
rect 30840 32376 30892 32385
rect 36452 32444 36504 32496
rect 36360 32419 36412 32428
rect 27804 32240 27856 32292
rect 31116 32308 31168 32360
rect 36360 32385 36369 32419
rect 36369 32385 36403 32419
rect 36403 32385 36412 32419
rect 36360 32376 36412 32385
rect 38660 32512 38712 32564
rect 39028 32512 39080 32564
rect 40040 32512 40092 32564
rect 40960 32512 41012 32564
rect 44824 32512 44876 32564
rect 38568 32419 38620 32428
rect 38568 32385 38577 32419
rect 38577 32385 38611 32419
rect 38611 32385 38620 32419
rect 38568 32376 38620 32385
rect 36176 32308 36228 32360
rect 36636 32351 36688 32360
rect 36636 32317 36645 32351
rect 36645 32317 36679 32351
rect 36679 32317 36688 32351
rect 37648 32351 37700 32360
rect 36636 32308 36688 32317
rect 37648 32317 37657 32351
rect 37657 32317 37691 32351
rect 37691 32317 37700 32351
rect 37648 32308 37700 32317
rect 38384 32351 38436 32360
rect 38384 32317 38393 32351
rect 38393 32317 38427 32351
rect 38427 32317 38436 32351
rect 38384 32308 38436 32317
rect 29184 32283 29236 32292
rect 29184 32249 29193 32283
rect 29193 32249 29227 32283
rect 29227 32249 29236 32283
rect 29184 32240 29236 32249
rect 30288 32240 30340 32292
rect 39764 32444 39816 32496
rect 39948 32376 40000 32428
rect 40316 32419 40368 32428
rect 40316 32385 40325 32419
rect 40325 32385 40359 32419
rect 40359 32385 40368 32419
rect 40316 32376 40368 32385
rect 41696 32376 41748 32428
rect 42432 32419 42484 32428
rect 42432 32385 42441 32419
rect 42441 32385 42475 32419
rect 42475 32385 42484 32419
rect 42432 32376 42484 32385
rect 43536 32419 43588 32428
rect 43536 32385 43545 32419
rect 43545 32385 43579 32419
rect 43579 32385 43588 32419
rect 43536 32376 43588 32385
rect 44456 32376 44508 32428
rect 47768 32419 47820 32428
rect 47768 32385 47777 32419
rect 47777 32385 47811 32419
rect 47811 32385 47820 32419
rect 47768 32376 47820 32385
rect 43352 32351 43404 32360
rect 43352 32317 43361 32351
rect 43361 32317 43395 32351
rect 43395 32317 43404 32351
rect 43352 32308 43404 32317
rect 24952 32172 25004 32224
rect 28632 32172 28684 32224
rect 32588 32172 32640 32224
rect 33876 32172 33928 32224
rect 46480 32240 46532 32292
rect 44180 32215 44232 32224
rect 44180 32181 44189 32215
rect 44189 32181 44223 32215
rect 44223 32181 44232 32215
rect 44180 32172 44232 32181
rect 47584 32215 47636 32224
rect 47584 32181 47593 32215
rect 47593 32181 47627 32215
rect 47627 32181 47636 32215
rect 47584 32172 47636 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2504 32011 2556 32020
rect 2504 31977 2513 32011
rect 2513 31977 2547 32011
rect 2547 31977 2556 32011
rect 2504 31968 2556 31977
rect 26056 32011 26108 32020
rect 26056 31977 26065 32011
rect 26065 31977 26099 32011
rect 26099 31977 26108 32011
rect 26056 31968 26108 31977
rect 29552 31968 29604 32020
rect 29276 31900 29328 31952
rect 24400 31832 24452 31884
rect 27620 31875 27672 31884
rect 27620 31841 27629 31875
rect 27629 31841 27663 31875
rect 27663 31841 27672 31875
rect 27620 31832 27672 31841
rect 8576 31764 8628 31816
rect 24952 31807 25004 31816
rect 24952 31773 24986 31807
rect 24986 31773 25004 31807
rect 24952 31764 25004 31773
rect 27804 31807 27856 31816
rect 27804 31773 27813 31807
rect 27813 31773 27847 31807
rect 27847 31773 27856 31807
rect 27804 31764 27856 31773
rect 28356 31764 28408 31816
rect 29184 31832 29236 31884
rect 29552 31875 29604 31884
rect 29552 31841 29561 31875
rect 29561 31841 29595 31875
rect 29595 31841 29604 31875
rect 29552 31832 29604 31841
rect 29000 31764 29052 31816
rect 29736 31764 29788 31816
rect 30104 31832 30156 31884
rect 31300 31764 31352 31816
rect 33048 31832 33100 31884
rect 35440 31968 35492 32020
rect 36176 32011 36228 32020
rect 36176 31977 36185 32011
rect 36185 31977 36219 32011
rect 36219 31977 36228 32011
rect 36176 31968 36228 31977
rect 36636 31968 36688 32020
rect 42800 32011 42852 32020
rect 42800 31977 42809 32011
rect 42809 31977 42843 32011
rect 42843 31977 42852 32011
rect 42800 31968 42852 31977
rect 43536 31968 43588 32020
rect 33784 31943 33836 31952
rect 33784 31909 33793 31943
rect 33793 31909 33827 31943
rect 33827 31909 33836 31943
rect 33784 31900 33836 31909
rect 28816 31739 28868 31748
rect 28816 31705 28825 31739
rect 28825 31705 28859 31739
rect 28859 31705 28868 31739
rect 28816 31696 28868 31705
rect 30104 31696 30156 31748
rect 32404 31807 32456 31816
rect 32404 31773 32413 31807
rect 32413 31773 32447 31807
rect 32447 31773 32456 31807
rect 32404 31764 32456 31773
rect 32588 31807 32640 31816
rect 32588 31773 32597 31807
rect 32597 31773 32631 31807
rect 32631 31773 32640 31807
rect 32588 31764 32640 31773
rect 32956 31764 33008 31816
rect 33140 31807 33192 31816
rect 33140 31773 33149 31807
rect 33149 31773 33183 31807
rect 33183 31773 33192 31807
rect 33140 31764 33192 31773
rect 34704 31832 34756 31884
rect 34428 31764 34480 31816
rect 37280 31900 37332 31952
rect 37648 31900 37700 31952
rect 38384 31900 38436 31952
rect 35900 31875 35952 31884
rect 35900 31841 35909 31875
rect 35909 31841 35943 31875
rect 35943 31841 35952 31875
rect 35900 31832 35952 31841
rect 37004 31832 37056 31884
rect 38016 31875 38068 31884
rect 34152 31696 34204 31748
rect 36544 31764 36596 31816
rect 37096 31807 37148 31816
rect 36912 31742 36964 31794
rect 37096 31773 37105 31807
rect 37105 31773 37139 31807
rect 37139 31773 37148 31807
rect 37096 31764 37148 31773
rect 38016 31841 38025 31875
rect 38025 31841 38059 31875
rect 38059 31841 38068 31875
rect 38016 31832 38068 31841
rect 38568 31764 38620 31816
rect 42524 31900 42576 31952
rect 39948 31875 40000 31884
rect 39948 31841 39957 31875
rect 39957 31841 39991 31875
rect 39991 31841 40000 31875
rect 39948 31832 40000 31841
rect 40408 31875 40460 31884
rect 40408 31841 40417 31875
rect 40417 31841 40451 31875
rect 40451 31841 40460 31875
rect 40408 31832 40460 31841
rect 41696 31832 41748 31884
rect 40040 31807 40092 31816
rect 40040 31773 40049 31807
rect 40049 31773 40083 31807
rect 40083 31773 40092 31807
rect 40040 31764 40092 31773
rect 41420 31807 41472 31816
rect 41420 31773 41429 31807
rect 41429 31773 41463 31807
rect 41463 31773 41472 31807
rect 42340 31807 42392 31816
rect 41420 31764 41472 31773
rect 42340 31773 42349 31807
rect 42349 31773 42383 31807
rect 42383 31773 42392 31807
rect 42340 31764 42392 31773
rect 43444 31764 43496 31816
rect 46940 31900 46992 31952
rect 46480 31875 46532 31884
rect 46480 31841 46489 31875
rect 46489 31841 46523 31875
rect 46523 31841 46532 31875
rect 46480 31832 46532 31841
rect 48136 31875 48188 31884
rect 48136 31841 48145 31875
rect 48145 31841 48179 31875
rect 48179 31841 48188 31875
rect 48136 31832 48188 31841
rect 40316 31696 40368 31748
rect 43628 31739 43680 31748
rect 43628 31705 43637 31739
rect 43637 31705 43671 31739
rect 43671 31705 43680 31739
rect 43628 31696 43680 31705
rect 27988 31671 28040 31680
rect 27988 31637 27997 31671
rect 27997 31637 28031 31671
rect 28031 31637 28040 31671
rect 27988 31628 28040 31637
rect 28908 31628 28960 31680
rect 32220 31628 32272 31680
rect 33968 31671 34020 31680
rect 33968 31637 33977 31671
rect 33977 31637 34011 31671
rect 34011 31637 34020 31671
rect 33968 31628 34020 31637
rect 37004 31671 37056 31680
rect 37004 31637 37013 31671
rect 37013 31637 37047 31671
rect 37047 31637 37056 31671
rect 37004 31628 37056 31637
rect 38844 31671 38896 31680
rect 38844 31637 38853 31671
rect 38853 31637 38887 31671
rect 38887 31637 38896 31671
rect 38844 31628 38896 31637
rect 41236 31671 41288 31680
rect 41236 31637 41245 31671
rect 41245 31637 41279 31671
rect 41279 31637 41288 31671
rect 41236 31628 41288 31637
rect 43168 31628 43220 31680
rect 43904 31671 43956 31680
rect 43904 31637 43913 31671
rect 43913 31637 43947 31671
rect 43947 31637 43956 31671
rect 43904 31628 43956 31637
rect 43996 31671 44048 31680
rect 43996 31637 44005 31671
rect 44005 31637 44039 31671
rect 44039 31637 44048 31671
rect 43996 31628 44048 31637
rect 44272 31628 44324 31680
rect 46940 31628 46992 31680
rect 48044 31628 48096 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 33784 31399 33836 31408
rect 23848 31331 23900 31340
rect 23848 31297 23857 31331
rect 23857 31297 23891 31331
rect 23891 31297 23900 31331
rect 23848 31288 23900 31297
rect 24216 31288 24268 31340
rect 24400 31288 24452 31340
rect 25136 31288 25188 31340
rect 29092 31288 29144 31340
rect 28908 31263 28960 31272
rect 28908 31229 28917 31263
rect 28917 31229 28951 31263
rect 28951 31229 28960 31263
rect 28908 31220 28960 31229
rect 29736 31288 29788 31340
rect 30104 31331 30156 31340
rect 30104 31297 30113 31331
rect 30113 31297 30147 31331
rect 30147 31297 30156 31331
rect 30288 31331 30340 31340
rect 30104 31288 30156 31297
rect 30288 31297 30297 31331
rect 30297 31297 30331 31331
rect 30331 31297 30340 31331
rect 30288 31288 30340 31297
rect 33784 31365 33818 31399
rect 33818 31365 33836 31399
rect 33784 31356 33836 31365
rect 31760 31288 31812 31340
rect 27988 31152 28040 31204
rect 28448 31152 28500 31204
rect 32036 31220 32088 31272
rect 34796 31424 34848 31476
rect 37004 31424 37056 31476
rect 42892 31424 42944 31476
rect 43352 31424 43404 31476
rect 43996 31424 44048 31476
rect 36176 31356 36228 31408
rect 36452 31356 36504 31408
rect 36912 31288 36964 31340
rect 40408 31356 40460 31408
rect 41236 31356 41288 31408
rect 38844 31331 38896 31340
rect 38844 31297 38853 31331
rect 38853 31297 38887 31331
rect 38887 31297 38896 31331
rect 39028 31331 39080 31340
rect 38844 31288 38896 31297
rect 39028 31297 39037 31331
rect 39037 31297 39071 31331
rect 39071 31297 39080 31331
rect 39028 31288 39080 31297
rect 41144 31288 41196 31340
rect 42892 31331 42944 31340
rect 42892 31297 42901 31331
rect 42901 31297 42935 31331
rect 42935 31297 42944 31331
rect 42892 31288 42944 31297
rect 43628 31356 43680 31408
rect 44180 31356 44232 31408
rect 47492 31424 47544 31476
rect 47768 31424 47820 31476
rect 46112 31356 46164 31408
rect 47032 31356 47084 31408
rect 43076 31263 43128 31272
rect 38752 31152 38804 31204
rect 43076 31229 43085 31263
rect 43085 31229 43119 31263
rect 43119 31229 43128 31263
rect 43904 31288 43956 31340
rect 45744 31331 45796 31340
rect 45744 31297 45753 31331
rect 45753 31297 45787 31331
rect 45787 31297 45796 31331
rect 45744 31288 45796 31297
rect 43812 31263 43864 31272
rect 43076 31220 43128 31229
rect 43812 31229 43821 31263
rect 43821 31229 43855 31263
rect 43855 31229 43864 31263
rect 43812 31220 43864 31229
rect 46020 31288 46072 31340
rect 46848 31288 46900 31340
rect 47308 31288 47360 31340
rect 48044 31220 48096 31272
rect 44824 31152 44876 31204
rect 24860 31084 24912 31136
rect 29276 31084 29328 31136
rect 29828 31127 29880 31136
rect 29828 31093 29837 31127
rect 29837 31093 29871 31127
rect 29871 31093 29880 31127
rect 29828 31084 29880 31093
rect 33508 31084 33560 31136
rect 34428 31084 34480 31136
rect 38844 31084 38896 31136
rect 41972 31084 42024 31136
rect 43168 31127 43220 31136
rect 43168 31093 43177 31127
rect 43177 31093 43211 31127
rect 43211 31093 43220 31127
rect 43168 31084 43220 31093
rect 45100 31084 45152 31136
rect 47768 31152 47820 31204
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 25136 30880 25188 30932
rect 28908 30880 28960 30932
rect 33968 30880 34020 30932
rect 34704 30923 34756 30932
rect 34704 30889 34713 30923
rect 34713 30889 34747 30923
rect 34747 30889 34756 30923
rect 34704 30880 34756 30889
rect 41420 30880 41472 30932
rect 42340 30923 42392 30932
rect 42340 30889 42349 30923
rect 42349 30889 42383 30923
rect 42383 30889 42392 30923
rect 42340 30880 42392 30889
rect 44456 30880 44508 30932
rect 46020 30923 46072 30932
rect 46020 30889 46029 30923
rect 46029 30889 46063 30923
rect 46063 30889 46072 30923
rect 46020 30880 46072 30889
rect 44180 30812 44232 30864
rect 47032 30880 47084 30932
rect 47492 30880 47544 30932
rect 33140 30744 33192 30796
rect 24860 30719 24912 30728
rect 24860 30685 24869 30719
rect 24869 30685 24903 30719
rect 24903 30685 24912 30719
rect 24860 30676 24912 30685
rect 28448 30719 28500 30728
rect 28448 30685 28457 30719
rect 28457 30685 28491 30719
rect 28491 30685 28500 30719
rect 28448 30676 28500 30685
rect 28816 30719 28868 30728
rect 28816 30685 28825 30719
rect 28825 30685 28859 30719
rect 28859 30685 28868 30719
rect 28816 30676 28868 30685
rect 32128 30719 32180 30728
rect 32128 30685 32137 30719
rect 32137 30685 32171 30719
rect 32171 30685 32180 30719
rect 32128 30676 32180 30685
rect 32220 30676 32272 30728
rect 34796 30676 34848 30728
rect 29000 30608 29052 30660
rect 27436 30540 27488 30592
rect 33508 30583 33560 30592
rect 33508 30549 33517 30583
rect 33517 30549 33551 30583
rect 33551 30549 33560 30583
rect 33508 30540 33560 30549
rect 39856 30744 39908 30796
rect 41604 30744 41656 30796
rect 41972 30787 42024 30796
rect 41972 30753 41981 30787
rect 41981 30753 42015 30787
rect 42015 30753 42024 30787
rect 41972 30744 42024 30753
rect 40132 30676 40184 30728
rect 41144 30719 41196 30728
rect 41144 30685 41153 30719
rect 41153 30685 41187 30719
rect 41187 30685 41196 30719
rect 41144 30676 41196 30685
rect 41420 30676 41472 30728
rect 42800 30744 42852 30796
rect 43076 30719 43128 30728
rect 43076 30685 43085 30719
rect 43085 30685 43119 30719
rect 43119 30685 43128 30719
rect 43076 30676 43128 30685
rect 44272 30744 44324 30796
rect 44364 30744 44416 30796
rect 44456 30719 44508 30728
rect 44456 30685 44465 30719
rect 44465 30685 44499 30719
rect 44499 30685 44508 30719
rect 44456 30676 44508 30685
rect 34980 30608 35032 30660
rect 37188 30608 37240 30660
rect 38108 30651 38160 30660
rect 38108 30617 38117 30651
rect 38117 30617 38151 30651
rect 38151 30617 38160 30651
rect 38108 30608 38160 30617
rect 39028 30608 39080 30660
rect 45652 30676 45704 30728
rect 46112 30719 46164 30728
rect 46112 30685 46121 30719
rect 46121 30685 46155 30719
rect 46155 30685 46164 30719
rect 46112 30676 46164 30685
rect 47584 30676 47636 30728
rect 36268 30540 36320 30592
rect 40408 30583 40460 30592
rect 40408 30549 40417 30583
rect 40417 30549 40451 30583
rect 40451 30549 40460 30583
rect 40408 30540 40460 30549
rect 40592 30540 40644 30592
rect 44824 30540 44876 30592
rect 45100 30608 45152 30660
rect 45744 30608 45796 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 30840 30268 30892 30320
rect 38936 30336 38988 30388
rect 41604 30336 41656 30388
rect 47032 30379 47084 30388
rect 47032 30345 47041 30379
rect 47041 30345 47075 30379
rect 47075 30345 47084 30379
rect 47032 30336 47084 30345
rect 29276 30243 29328 30252
rect 29276 30209 29285 30243
rect 29285 30209 29319 30243
rect 29319 30209 29328 30243
rect 29276 30200 29328 30209
rect 29460 30243 29512 30252
rect 29460 30209 29469 30243
rect 29469 30209 29503 30243
rect 29503 30209 29512 30243
rect 29460 30200 29512 30209
rect 35440 30200 35492 30252
rect 40408 30268 40460 30320
rect 41420 30311 41472 30320
rect 41420 30277 41429 30311
rect 41429 30277 41463 30311
rect 41463 30277 41472 30311
rect 41420 30268 41472 30277
rect 36544 30243 36596 30252
rect 36544 30209 36553 30243
rect 36553 30209 36587 30243
rect 36587 30209 36596 30243
rect 36544 30200 36596 30209
rect 36728 30243 36780 30252
rect 36728 30209 36737 30243
rect 36737 30209 36771 30243
rect 36771 30209 36780 30243
rect 37280 30243 37332 30252
rect 36728 30200 36780 30209
rect 37280 30209 37289 30243
rect 37289 30209 37323 30243
rect 37323 30209 37332 30243
rect 37280 30200 37332 30209
rect 37372 30200 37424 30252
rect 37556 30243 37608 30252
rect 37556 30209 37565 30243
rect 37565 30209 37599 30243
rect 37599 30209 37608 30243
rect 37556 30200 37608 30209
rect 38568 30200 38620 30252
rect 38752 30243 38804 30252
rect 38752 30209 38761 30243
rect 38761 30209 38795 30243
rect 38795 30209 38804 30243
rect 38752 30200 38804 30209
rect 38844 30200 38896 30252
rect 43812 30268 43864 30320
rect 42524 30200 42576 30252
rect 47768 30243 47820 30252
rect 33416 30064 33468 30116
rect 43812 30132 43864 30184
rect 45652 30175 45704 30184
rect 45652 30141 45661 30175
rect 45661 30141 45695 30175
rect 45695 30141 45704 30175
rect 45652 30132 45704 30141
rect 37648 30064 37700 30116
rect 40316 30064 40368 30116
rect 41604 30107 41656 30116
rect 41604 30073 41613 30107
rect 41613 30073 41647 30107
rect 41647 30073 41656 30107
rect 41604 30064 41656 30073
rect 47768 30209 47777 30243
rect 47777 30209 47811 30243
rect 47811 30209 47820 30243
rect 47768 30200 47820 30209
rect 30012 29996 30064 30048
rect 36084 30039 36136 30048
rect 36084 30005 36093 30039
rect 36093 30005 36127 30039
rect 36127 30005 36136 30039
rect 36084 29996 36136 30005
rect 37832 30039 37884 30048
rect 37832 30005 37841 30039
rect 37841 30005 37875 30039
rect 37875 30005 37884 30039
rect 37832 29996 37884 30005
rect 43904 29996 43956 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 36820 29792 36872 29844
rect 38936 29792 38988 29844
rect 40500 29835 40552 29844
rect 40500 29801 40509 29835
rect 40509 29801 40543 29835
rect 40543 29801 40552 29835
rect 40500 29792 40552 29801
rect 43444 29835 43496 29844
rect 43444 29801 43453 29835
rect 43453 29801 43487 29835
rect 43487 29801 43496 29835
rect 43444 29792 43496 29801
rect 35900 29724 35952 29776
rect 22652 29588 22704 29640
rect 24676 29631 24728 29640
rect 24676 29597 24685 29631
rect 24685 29597 24719 29631
rect 24719 29597 24728 29631
rect 24676 29588 24728 29597
rect 24860 29631 24912 29640
rect 24860 29597 24874 29631
rect 24874 29597 24908 29631
rect 24908 29597 24912 29631
rect 24860 29588 24912 29597
rect 25596 29631 25648 29640
rect 25596 29597 25605 29631
rect 25605 29597 25639 29631
rect 25639 29597 25648 29631
rect 25596 29588 25648 29597
rect 26332 29588 26384 29640
rect 29276 29656 29328 29708
rect 30012 29699 30064 29708
rect 30012 29665 30021 29699
rect 30021 29665 30055 29699
rect 30055 29665 30064 29699
rect 30012 29656 30064 29665
rect 32956 29656 33008 29708
rect 37556 29656 37608 29708
rect 38016 29656 38068 29708
rect 29828 29588 29880 29640
rect 24400 29495 24452 29504
rect 24400 29461 24409 29495
rect 24409 29461 24443 29495
rect 24443 29461 24452 29495
rect 24400 29452 24452 29461
rect 24768 29452 24820 29504
rect 24860 29452 24912 29504
rect 25872 29563 25924 29572
rect 25872 29529 25906 29563
rect 25906 29529 25924 29563
rect 25872 29520 25924 29529
rect 32128 29588 32180 29640
rect 33416 29631 33468 29640
rect 25964 29452 26016 29504
rect 28816 29452 28868 29504
rect 30932 29452 30984 29504
rect 31484 29452 31536 29504
rect 32128 29452 32180 29504
rect 33416 29597 33425 29631
rect 33425 29597 33459 29631
rect 33459 29597 33468 29631
rect 33416 29588 33468 29597
rect 33508 29588 33560 29640
rect 34336 29588 34388 29640
rect 34704 29588 34756 29640
rect 35348 29588 35400 29640
rect 36084 29588 36136 29640
rect 37372 29588 37424 29640
rect 38568 29631 38620 29640
rect 38568 29597 38577 29631
rect 38577 29597 38611 29631
rect 38611 29597 38620 29631
rect 38568 29588 38620 29597
rect 40316 29724 40368 29776
rect 33784 29520 33836 29572
rect 34152 29563 34204 29572
rect 34152 29529 34161 29563
rect 34161 29529 34195 29563
rect 34195 29529 34204 29563
rect 34152 29520 34204 29529
rect 41144 29588 41196 29640
rect 43444 29588 43496 29640
rect 46296 29631 46348 29640
rect 46296 29597 46305 29631
rect 46305 29597 46339 29631
rect 46339 29597 46348 29631
rect 46296 29588 46348 29597
rect 40132 29563 40184 29572
rect 40132 29529 40141 29563
rect 40141 29529 40175 29563
rect 40175 29529 40184 29563
rect 40132 29520 40184 29529
rect 40224 29563 40276 29572
rect 40224 29529 40233 29563
rect 40233 29529 40267 29563
rect 40267 29529 40276 29563
rect 40224 29520 40276 29529
rect 43260 29520 43312 29572
rect 46480 29563 46532 29572
rect 46480 29529 46489 29563
rect 46489 29529 46523 29563
rect 46523 29529 46532 29563
rect 46480 29520 46532 29529
rect 48136 29563 48188 29572
rect 48136 29529 48145 29563
rect 48145 29529 48179 29563
rect 48179 29529 48188 29563
rect 48136 29520 48188 29529
rect 33140 29452 33192 29504
rect 33232 29452 33284 29504
rect 33600 29452 33652 29504
rect 37280 29452 37332 29504
rect 37924 29452 37976 29504
rect 44272 29452 44324 29504
rect 44456 29452 44508 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 18880 29248 18932 29300
rect 24584 29248 24636 29300
rect 24676 29248 24728 29300
rect 25872 29248 25924 29300
rect 26240 29248 26292 29300
rect 27620 29248 27672 29300
rect 17776 29155 17828 29164
rect 17776 29121 17785 29155
rect 17785 29121 17819 29155
rect 17819 29121 17828 29155
rect 17776 29112 17828 29121
rect 23204 29112 23256 29164
rect 24860 29180 24912 29232
rect 24400 29112 24452 29164
rect 25872 29112 25924 29164
rect 29460 29248 29512 29300
rect 33232 29248 33284 29300
rect 35348 29291 35400 29300
rect 22652 29087 22704 29096
rect 22652 29053 22661 29087
rect 22661 29053 22695 29087
rect 22695 29053 22704 29087
rect 22652 29044 22704 29053
rect 25780 29044 25832 29096
rect 26332 29155 26384 29164
rect 26332 29121 26341 29155
rect 26341 29121 26375 29155
rect 26375 29121 26384 29155
rect 27436 29155 27488 29164
rect 26332 29112 26384 29121
rect 27436 29121 27445 29155
rect 27445 29121 27479 29155
rect 27479 29121 27488 29155
rect 27436 29112 27488 29121
rect 28080 29155 28132 29164
rect 28080 29121 28089 29155
rect 28089 29121 28123 29155
rect 28123 29121 28132 29155
rect 28080 29112 28132 29121
rect 28172 29112 28224 29164
rect 29920 29155 29972 29164
rect 29920 29121 29929 29155
rect 29929 29121 29963 29155
rect 29963 29121 29972 29155
rect 29920 29112 29972 29121
rect 32128 29180 32180 29232
rect 33600 29180 33652 29232
rect 30932 29155 30984 29164
rect 30932 29121 30941 29155
rect 30941 29121 30975 29155
rect 30975 29121 30984 29155
rect 30932 29112 30984 29121
rect 31760 29112 31812 29164
rect 33692 29112 33744 29164
rect 34428 29180 34480 29232
rect 35348 29257 35357 29291
rect 35357 29257 35391 29291
rect 35391 29257 35400 29291
rect 35348 29248 35400 29257
rect 41144 29291 41196 29300
rect 41144 29257 41153 29291
rect 41153 29257 41187 29291
rect 41187 29257 41196 29291
rect 41144 29248 41196 29257
rect 43444 29291 43496 29300
rect 43444 29257 43453 29291
rect 43453 29257 43487 29291
rect 43487 29257 43496 29291
rect 43444 29248 43496 29257
rect 34336 29155 34388 29164
rect 34336 29121 34361 29155
rect 34361 29121 34388 29155
rect 23480 28976 23532 29028
rect 26056 28976 26108 29028
rect 22928 28908 22980 28960
rect 26700 28908 26752 28960
rect 27528 28951 27580 28960
rect 27528 28917 27537 28951
rect 27537 28917 27571 28951
rect 27571 28917 27580 28951
rect 27528 28908 27580 28917
rect 33508 29044 33560 29096
rect 28724 28908 28776 28960
rect 29460 28951 29512 28960
rect 29460 28917 29469 28951
rect 29469 28917 29503 28951
rect 29503 28917 29512 28951
rect 29460 28908 29512 28917
rect 34336 29112 34388 29121
rect 34796 29155 34848 29164
rect 34796 29121 34805 29155
rect 34805 29121 34839 29155
rect 34839 29121 34848 29155
rect 34796 29112 34848 29121
rect 35900 29180 35952 29232
rect 37004 29180 37056 29232
rect 45008 29248 45060 29300
rect 44180 29223 44232 29232
rect 36360 29155 36412 29164
rect 34428 29044 34480 29096
rect 36360 29121 36369 29155
rect 36369 29121 36403 29155
rect 36403 29121 36412 29155
rect 36360 29112 36412 29121
rect 37280 29155 37332 29164
rect 35992 29044 36044 29096
rect 37280 29121 37289 29155
rect 37289 29121 37323 29155
rect 37323 29121 37332 29155
rect 37280 29112 37332 29121
rect 37648 29112 37700 29164
rect 40592 29112 40644 29164
rect 44180 29189 44214 29223
rect 44214 29189 44232 29223
rect 44180 29180 44232 29189
rect 43352 29112 43404 29164
rect 46296 29112 46348 29164
rect 37464 29044 37516 29096
rect 43812 29044 43864 29096
rect 34244 29019 34296 29028
rect 34244 28985 34253 29019
rect 34253 28985 34287 29019
rect 34287 28985 34296 29019
rect 34244 28976 34296 28985
rect 40500 28976 40552 29028
rect 40776 28976 40828 29028
rect 34428 28908 34480 28960
rect 36176 28951 36228 28960
rect 36176 28917 36185 28951
rect 36185 28917 36219 28951
rect 36219 28917 36228 28951
rect 36176 28908 36228 28917
rect 40224 28951 40276 28960
rect 40224 28917 40233 28951
rect 40233 28917 40267 28951
rect 40267 28917 40276 28951
rect 40224 28908 40276 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19984 28747 20036 28756
rect 19984 28713 19993 28747
rect 19993 28713 20027 28747
rect 20027 28713 20036 28747
rect 19984 28704 20036 28713
rect 24952 28704 25004 28756
rect 26148 28704 26200 28756
rect 26240 28704 26292 28756
rect 26700 28704 26752 28756
rect 18512 28611 18564 28620
rect 18512 28577 18521 28611
rect 18521 28577 18555 28611
rect 18555 28577 18564 28611
rect 18512 28568 18564 28577
rect 18788 28568 18840 28620
rect 22652 28500 22704 28552
rect 22836 28543 22888 28552
rect 22836 28509 22845 28543
rect 22845 28509 22879 28543
rect 22879 28509 22888 28543
rect 22836 28500 22888 28509
rect 17132 28475 17184 28484
rect 17132 28441 17141 28475
rect 17141 28441 17175 28475
rect 17175 28441 17184 28475
rect 17132 28432 17184 28441
rect 17776 28475 17828 28484
rect 17776 28441 17785 28475
rect 17785 28441 17819 28475
rect 17819 28441 17828 28475
rect 17776 28432 17828 28441
rect 24768 28636 24820 28688
rect 28172 28704 28224 28756
rect 34796 28704 34848 28756
rect 37372 28704 37424 28756
rect 37464 28704 37516 28756
rect 38568 28704 38620 28756
rect 40132 28704 40184 28756
rect 44088 28704 44140 28756
rect 44548 28704 44600 28756
rect 23756 28432 23808 28484
rect 22100 28407 22152 28416
rect 22100 28373 22109 28407
rect 22109 28373 22143 28407
rect 22143 28373 22152 28407
rect 22100 28364 22152 28373
rect 26148 28568 26200 28620
rect 25320 28500 25372 28552
rect 26056 28500 26108 28552
rect 26332 28543 26384 28552
rect 26332 28509 26341 28543
rect 26341 28509 26375 28543
rect 26375 28509 26384 28543
rect 26332 28500 26384 28509
rect 27436 28543 27488 28552
rect 27436 28509 27445 28543
rect 27445 28509 27479 28543
rect 27479 28509 27488 28543
rect 27436 28500 27488 28509
rect 33692 28636 33744 28688
rect 34704 28636 34756 28688
rect 29460 28568 29512 28620
rect 33508 28568 33560 28620
rect 40500 28636 40552 28688
rect 28540 28543 28592 28552
rect 28540 28509 28549 28543
rect 28549 28509 28583 28543
rect 28583 28509 28592 28543
rect 28540 28500 28592 28509
rect 28724 28543 28776 28552
rect 28724 28509 28733 28543
rect 28733 28509 28767 28543
rect 28767 28509 28776 28543
rect 33876 28543 33928 28552
rect 28724 28500 28776 28509
rect 33876 28509 33885 28543
rect 33885 28509 33919 28543
rect 33919 28509 33928 28543
rect 33876 28500 33928 28509
rect 35900 28500 35952 28552
rect 36360 28500 36412 28552
rect 37832 28568 37884 28620
rect 44732 28568 44784 28620
rect 47676 28568 47728 28620
rect 37004 28500 37056 28552
rect 37648 28543 37700 28552
rect 37648 28509 37657 28543
rect 37657 28509 37691 28543
rect 37691 28509 37700 28543
rect 37648 28500 37700 28509
rect 38108 28500 38160 28552
rect 40040 28500 40092 28552
rect 40684 28500 40736 28552
rect 40868 28500 40920 28552
rect 43352 28543 43404 28552
rect 43352 28509 43361 28543
rect 43361 28509 43395 28543
rect 43395 28509 43404 28543
rect 43352 28500 43404 28509
rect 33140 28432 33192 28484
rect 34152 28432 34204 28484
rect 34244 28432 34296 28484
rect 35992 28432 36044 28484
rect 36176 28432 36228 28484
rect 42984 28432 43036 28484
rect 46940 28432 46992 28484
rect 48136 28475 48188 28484
rect 48136 28441 48145 28475
rect 48145 28441 48179 28475
rect 48179 28441 48188 28475
rect 48136 28432 48188 28441
rect 27620 28364 27672 28416
rect 29552 28364 29604 28416
rect 34612 28364 34664 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 16764 28160 16816 28212
rect 17132 28160 17184 28212
rect 22836 28203 22888 28212
rect 18144 28135 18196 28144
rect 18144 28101 18153 28135
rect 18153 28101 18187 28135
rect 18187 28101 18196 28135
rect 18144 28092 18196 28101
rect 18420 28092 18472 28144
rect 22836 28169 22845 28203
rect 22845 28169 22879 28203
rect 22879 28169 22888 28203
rect 22836 28160 22888 28169
rect 26332 28160 26384 28212
rect 27436 28160 27488 28212
rect 28540 28160 28592 28212
rect 31760 28160 31812 28212
rect 32404 28160 32456 28212
rect 34428 28160 34480 28212
rect 35900 28160 35952 28212
rect 40592 28203 40644 28212
rect 40592 28169 40601 28203
rect 40601 28169 40635 28203
rect 40635 28169 40644 28203
rect 40592 28160 40644 28169
rect 41236 28160 41288 28212
rect 46480 28160 46532 28212
rect 31944 28092 31996 28144
rect 32312 28135 32364 28144
rect 32312 28101 32321 28135
rect 32321 28101 32355 28135
rect 32355 28101 32364 28135
rect 32312 28092 32364 28101
rect 17040 28067 17092 28076
rect 17040 28033 17049 28067
rect 17049 28033 17083 28067
rect 17083 28033 17092 28067
rect 17040 28024 17092 28033
rect 17776 28067 17828 28076
rect 17776 28033 17785 28067
rect 17785 28033 17819 28067
rect 17819 28033 17828 28067
rect 17776 28024 17828 28033
rect 22100 28024 22152 28076
rect 23480 28067 23532 28076
rect 23480 28033 23489 28067
rect 23489 28033 23523 28067
rect 23523 28033 23532 28067
rect 23480 28024 23532 28033
rect 23756 28067 23808 28076
rect 23756 28033 23765 28067
rect 23765 28033 23799 28067
rect 23799 28033 23808 28067
rect 23756 28024 23808 28033
rect 26148 28024 26200 28076
rect 26424 28024 26476 28076
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 29368 28024 29420 28076
rect 30380 28024 30432 28076
rect 22560 27999 22612 28008
rect 22560 27965 22569 27999
rect 22569 27965 22603 27999
rect 22603 27965 22612 27999
rect 22560 27956 22612 27965
rect 25964 27999 26016 28008
rect 25964 27965 25973 27999
rect 25973 27965 26007 27999
rect 26007 27965 26016 27999
rect 25964 27956 26016 27965
rect 28724 27999 28776 28008
rect 25228 27888 25280 27940
rect 28724 27965 28733 27999
rect 28733 27965 28767 27999
rect 28767 27965 28776 27999
rect 28724 27956 28776 27965
rect 27988 27888 28040 27940
rect 29920 27888 29972 27940
rect 31484 28024 31536 28076
rect 31852 28024 31904 28076
rect 32404 28067 32456 28076
rect 32404 28033 32413 28067
rect 32413 28033 32447 28067
rect 32447 28033 32456 28067
rect 33876 28067 33928 28076
rect 32404 28024 32456 28033
rect 33876 28033 33885 28067
rect 33885 28033 33919 28067
rect 33919 28033 33928 28067
rect 33876 28024 33928 28033
rect 34704 28024 34756 28076
rect 40224 28024 40276 28076
rect 40776 28024 40828 28076
rect 41144 28067 41196 28076
rect 41144 28033 41153 28067
rect 41153 28033 41187 28067
rect 41187 28033 41196 28067
rect 41144 28024 41196 28033
rect 44272 28092 44324 28144
rect 36636 27956 36688 28008
rect 42432 27956 42484 28008
rect 42616 27956 42668 28008
rect 33324 27888 33376 27940
rect 33692 27888 33744 27940
rect 45836 28024 45888 28076
rect 46388 28067 46440 28076
rect 46388 28033 46397 28067
rect 46397 28033 46431 28067
rect 46431 28033 46440 28067
rect 46388 28024 46440 28033
rect 22652 27820 22704 27872
rect 24952 27820 25004 27872
rect 29552 27863 29604 27872
rect 29552 27829 29561 27863
rect 29561 27829 29595 27863
rect 29595 27829 29604 27863
rect 29552 27820 29604 27829
rect 31116 27863 31168 27872
rect 31116 27829 31125 27863
rect 31125 27829 31159 27863
rect 31159 27829 31168 27863
rect 31116 27820 31168 27829
rect 33140 27820 33192 27872
rect 40592 27820 40644 27872
rect 41512 27820 41564 27872
rect 43812 27820 43864 27872
rect 45284 27820 45336 27872
rect 46480 27863 46532 27872
rect 46480 27829 46489 27863
rect 46489 27829 46523 27863
rect 46523 27829 46532 27863
rect 46480 27820 46532 27829
rect 47768 27863 47820 27872
rect 47768 27829 47777 27863
rect 47777 27829 47811 27863
rect 47811 27829 47820 27863
rect 47768 27820 47820 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 26148 27659 26200 27668
rect 26148 27625 26157 27659
rect 26157 27625 26191 27659
rect 26191 27625 26200 27659
rect 26148 27616 26200 27625
rect 28724 27616 28776 27668
rect 34244 27616 34296 27668
rect 37648 27616 37700 27668
rect 23756 27548 23808 27600
rect 26056 27548 26108 27600
rect 26424 27548 26476 27600
rect 26516 27548 26568 27600
rect 25504 27480 25556 27532
rect 29368 27548 29420 27600
rect 34612 27548 34664 27600
rect 8392 27412 8444 27464
rect 17040 27412 17092 27464
rect 18052 27455 18104 27464
rect 18052 27421 18061 27455
rect 18061 27421 18095 27455
rect 18095 27421 18104 27455
rect 18052 27412 18104 27421
rect 25136 27455 25188 27464
rect 25136 27421 25145 27455
rect 25145 27421 25179 27455
rect 25179 27421 25188 27455
rect 25136 27412 25188 27421
rect 25596 27412 25648 27464
rect 26056 27455 26108 27464
rect 26056 27421 26065 27455
rect 26065 27421 26099 27455
rect 26099 27421 26108 27455
rect 26056 27412 26108 27421
rect 17316 27387 17368 27396
rect 17316 27353 17325 27387
rect 17325 27353 17359 27387
rect 17359 27353 17368 27387
rect 17316 27344 17368 27353
rect 18604 27387 18656 27396
rect 18604 27353 18613 27387
rect 18613 27353 18647 27387
rect 18647 27353 18656 27387
rect 18604 27344 18656 27353
rect 24124 27344 24176 27396
rect 25504 27276 25556 27328
rect 27160 27412 27212 27464
rect 28632 27344 28684 27396
rect 28908 27412 28960 27464
rect 28908 27276 28960 27328
rect 34428 27480 34480 27532
rect 37372 27523 37424 27532
rect 37372 27489 37381 27523
rect 37381 27489 37415 27523
rect 37415 27489 37424 27523
rect 37372 27480 37424 27489
rect 37648 27480 37700 27532
rect 32956 27412 33008 27464
rect 33692 27412 33744 27464
rect 34704 27455 34756 27464
rect 34704 27421 34713 27455
rect 34713 27421 34747 27455
rect 34747 27421 34756 27455
rect 34704 27412 34756 27421
rect 31116 27387 31168 27396
rect 31116 27353 31150 27387
rect 31150 27353 31168 27387
rect 31116 27344 31168 27353
rect 34888 27344 34940 27396
rect 35624 27455 35676 27464
rect 35624 27421 35633 27455
rect 35633 27421 35667 27455
rect 35667 27421 35676 27455
rect 35624 27412 35676 27421
rect 37280 27412 37332 27464
rect 38568 27548 38620 27600
rect 41144 27616 41196 27668
rect 39488 27548 39540 27600
rect 39212 27480 39264 27532
rect 39396 27480 39448 27532
rect 38108 27387 38160 27396
rect 31852 27276 31904 27328
rect 32220 27319 32272 27328
rect 32220 27285 32229 27319
rect 32229 27285 32263 27319
rect 32263 27285 32272 27319
rect 32220 27276 32272 27285
rect 33140 27276 33192 27328
rect 38108 27353 38117 27387
rect 38117 27353 38151 27387
rect 38151 27353 38160 27387
rect 38108 27344 38160 27353
rect 39488 27412 39540 27464
rect 47768 27548 47820 27600
rect 46480 27523 46532 27532
rect 46480 27489 46489 27523
rect 46489 27489 46523 27523
rect 46523 27489 46532 27523
rect 46480 27480 46532 27489
rect 46848 27523 46900 27532
rect 46848 27489 46857 27523
rect 46857 27489 46891 27523
rect 46891 27489 46900 27523
rect 46848 27480 46900 27489
rect 40316 27344 40368 27396
rect 43812 27412 43864 27464
rect 40868 27344 40920 27396
rect 35532 27319 35584 27328
rect 35532 27285 35541 27319
rect 35541 27285 35575 27319
rect 35575 27285 35584 27319
rect 35532 27276 35584 27285
rect 37004 27319 37056 27328
rect 37004 27285 37013 27319
rect 37013 27285 37047 27319
rect 37047 27285 37056 27319
rect 37004 27276 37056 27285
rect 37372 27276 37424 27328
rect 38476 27276 38528 27328
rect 38568 27276 38620 27328
rect 40776 27276 40828 27328
rect 41512 27344 41564 27396
rect 42892 27344 42944 27396
rect 46020 27344 46072 27396
rect 43444 27319 43496 27328
rect 43444 27285 43453 27319
rect 43453 27285 43487 27319
rect 43487 27285 43496 27319
rect 43444 27276 43496 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 16948 27072 17000 27124
rect 17040 27072 17092 27124
rect 8392 27004 8444 27056
rect 21916 27004 21968 27056
rect 25412 27004 25464 27056
rect 16672 26936 16724 26988
rect 18052 26979 18104 26988
rect 18052 26945 18061 26979
rect 18061 26945 18095 26979
rect 18095 26945 18104 26979
rect 18052 26936 18104 26945
rect 17868 26868 17920 26920
rect 22560 26868 22612 26920
rect 23020 26868 23072 26920
rect 7932 26775 7984 26784
rect 7932 26741 7941 26775
rect 7941 26741 7975 26775
rect 7975 26741 7984 26775
rect 7932 26732 7984 26741
rect 25136 26936 25188 26988
rect 26792 26936 26844 26988
rect 28264 26936 28316 26988
rect 28632 26979 28684 26988
rect 28632 26945 28641 26979
rect 28641 26945 28675 26979
rect 28675 26945 28684 26979
rect 28632 26936 28684 26945
rect 28908 26936 28960 26988
rect 24952 26868 25004 26920
rect 25780 26868 25832 26920
rect 25136 26843 25188 26852
rect 25136 26809 25145 26843
rect 25145 26809 25179 26843
rect 25179 26809 25188 26843
rect 25136 26800 25188 26809
rect 26424 26843 26476 26852
rect 26424 26809 26433 26843
rect 26433 26809 26467 26843
rect 26467 26809 26476 26843
rect 26424 26800 26476 26809
rect 27160 26868 27212 26920
rect 28540 26911 28592 26920
rect 28540 26877 28549 26911
rect 28549 26877 28583 26911
rect 28583 26877 28592 26911
rect 28540 26868 28592 26877
rect 32956 26936 33008 26988
rect 35532 27004 35584 27056
rect 37648 27004 37700 27056
rect 43352 27072 43404 27124
rect 46940 27115 46992 27124
rect 46940 27081 46949 27115
rect 46949 27081 46983 27115
rect 46983 27081 46992 27115
rect 46940 27072 46992 27081
rect 44088 27047 44140 27056
rect 28448 26800 28500 26852
rect 32680 26800 32732 26852
rect 27068 26732 27120 26784
rect 32864 26775 32916 26784
rect 32864 26741 32873 26775
rect 32873 26741 32907 26775
rect 32907 26741 32916 26775
rect 32864 26732 32916 26741
rect 33140 26911 33192 26920
rect 33140 26877 33149 26911
rect 33149 26877 33183 26911
rect 33183 26877 33192 26911
rect 36544 26936 36596 26988
rect 37372 26936 37424 26988
rect 37832 26936 37884 26988
rect 38568 26936 38620 26988
rect 38752 26936 38804 26988
rect 39856 26979 39908 26988
rect 39856 26945 39865 26979
rect 39865 26945 39899 26979
rect 39899 26945 39908 26979
rect 39856 26936 39908 26945
rect 40408 26936 40460 26988
rect 40684 26936 40736 26988
rect 41604 26936 41656 26988
rect 42892 26936 42944 26988
rect 44088 27013 44122 27047
rect 44122 27013 44140 27047
rect 44088 27004 44140 27013
rect 46112 26936 46164 26988
rect 33140 26868 33192 26877
rect 37648 26868 37700 26920
rect 43812 26911 43864 26920
rect 43812 26877 43821 26911
rect 43821 26877 43855 26911
rect 43855 26877 43864 26911
rect 43812 26868 43864 26877
rect 45376 26868 45428 26920
rect 47584 26936 47636 26988
rect 47676 26936 47728 26988
rect 35164 26800 35216 26852
rect 37280 26843 37332 26852
rect 34428 26732 34480 26784
rect 34796 26732 34848 26784
rect 37280 26809 37289 26843
rect 37289 26809 37323 26843
rect 37323 26809 37332 26843
rect 37280 26800 37332 26809
rect 41236 26843 41288 26852
rect 41236 26809 41245 26843
rect 41245 26809 41279 26843
rect 41279 26809 41288 26843
rect 41236 26800 41288 26809
rect 38016 26732 38068 26784
rect 38200 26732 38252 26784
rect 45744 26732 45796 26784
rect 46296 26732 46348 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8208 26528 8260 26580
rect 25412 26528 25464 26580
rect 25596 26571 25648 26580
rect 25596 26537 25605 26571
rect 25605 26537 25639 26571
rect 25639 26537 25648 26571
rect 25596 26528 25648 26537
rect 25964 26571 26016 26580
rect 25964 26537 25973 26571
rect 25973 26537 26007 26571
rect 26007 26537 26016 26571
rect 25964 26528 26016 26537
rect 26792 26571 26844 26580
rect 26792 26537 26801 26571
rect 26801 26537 26835 26571
rect 26835 26537 26844 26571
rect 26792 26528 26844 26537
rect 28632 26528 28684 26580
rect 40408 26571 40460 26580
rect 8208 26435 8260 26444
rect 8208 26401 8217 26435
rect 8217 26401 8251 26435
rect 8251 26401 8260 26435
rect 8208 26392 8260 26401
rect 17040 26392 17092 26444
rect 7932 26324 7984 26376
rect 16672 26367 16724 26376
rect 16672 26333 16681 26367
rect 16681 26333 16715 26367
rect 16715 26333 16724 26367
rect 16672 26324 16724 26333
rect 17316 26256 17368 26308
rect 33416 26460 33468 26512
rect 33692 26503 33744 26512
rect 33692 26469 33701 26503
rect 33701 26469 33735 26503
rect 33735 26469 33744 26503
rect 33692 26460 33744 26469
rect 35624 26460 35676 26512
rect 36268 26460 36320 26512
rect 37740 26460 37792 26512
rect 38292 26503 38344 26512
rect 38292 26469 38301 26503
rect 38301 26469 38335 26503
rect 38335 26469 38344 26503
rect 38292 26460 38344 26469
rect 40408 26537 40417 26571
rect 40417 26537 40451 26571
rect 40451 26537 40460 26571
rect 40408 26528 40460 26537
rect 40776 26571 40828 26580
rect 40776 26537 40785 26571
rect 40785 26537 40819 26571
rect 40819 26537 40828 26571
rect 40776 26528 40828 26537
rect 45376 26528 45428 26580
rect 45560 26528 45612 26580
rect 45928 26528 45980 26580
rect 23204 26435 23256 26444
rect 23204 26401 23213 26435
rect 23213 26401 23247 26435
rect 23247 26401 23256 26435
rect 23204 26392 23256 26401
rect 25228 26392 25280 26444
rect 25964 26392 26016 26444
rect 28356 26435 28408 26444
rect 23020 26367 23072 26376
rect 23020 26333 23029 26367
rect 23029 26333 23063 26367
rect 23063 26333 23072 26367
rect 25780 26367 25832 26376
rect 23020 26324 23072 26333
rect 25780 26333 25789 26367
rect 25789 26333 25823 26367
rect 25823 26333 25832 26367
rect 25780 26324 25832 26333
rect 26240 26324 26292 26376
rect 28356 26401 28365 26435
rect 28365 26401 28399 26435
rect 28399 26401 28408 26435
rect 28356 26392 28408 26401
rect 34704 26435 34756 26444
rect 34704 26401 34713 26435
rect 34713 26401 34747 26435
rect 34747 26401 34756 26435
rect 34704 26392 34756 26401
rect 37648 26392 37700 26444
rect 29644 26324 29696 26376
rect 32312 26367 32364 26376
rect 32312 26333 32321 26367
rect 32321 26333 32355 26367
rect 32355 26333 32364 26367
rect 32312 26324 32364 26333
rect 32956 26324 33008 26376
rect 34428 26324 34480 26376
rect 37832 26324 37884 26376
rect 32864 26256 32916 26308
rect 37004 26256 37056 26308
rect 37740 26256 37792 26308
rect 28172 26188 28224 26240
rect 29460 26188 29512 26240
rect 29736 26188 29788 26240
rect 33140 26188 33192 26240
rect 36452 26188 36504 26240
rect 38108 26256 38160 26308
rect 41236 26392 41288 26444
rect 45836 26460 45888 26512
rect 46940 26460 46992 26512
rect 38568 26367 38620 26376
rect 38568 26333 38577 26367
rect 38577 26333 38611 26367
rect 38611 26333 38620 26367
rect 38568 26324 38620 26333
rect 39948 26324 40000 26376
rect 40224 26324 40276 26376
rect 40592 26367 40644 26376
rect 40592 26333 40601 26367
rect 40601 26333 40635 26367
rect 40635 26333 40644 26367
rect 40592 26324 40644 26333
rect 43812 26392 43864 26444
rect 45652 26392 45704 26444
rect 46296 26435 46348 26444
rect 46296 26401 46305 26435
rect 46305 26401 46339 26435
rect 46339 26401 46348 26435
rect 46296 26392 46348 26401
rect 45008 26367 45060 26376
rect 45008 26333 45017 26367
rect 45017 26333 45051 26367
rect 45051 26333 45060 26367
rect 45008 26324 45060 26333
rect 45284 26367 45336 26376
rect 45284 26333 45293 26367
rect 45293 26333 45327 26367
rect 45327 26333 45336 26367
rect 45284 26324 45336 26333
rect 45744 26324 45796 26376
rect 45928 26324 45980 26376
rect 41604 26299 41656 26308
rect 41604 26265 41613 26299
rect 41613 26265 41647 26299
rect 41647 26265 41656 26299
rect 41604 26256 41656 26265
rect 44732 26256 44784 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 26240 26027 26292 26036
rect 26240 25993 26249 26027
rect 26249 25993 26283 26027
rect 26283 25993 26292 26027
rect 26240 25984 26292 25993
rect 27068 26027 27120 26036
rect 27068 25993 27077 26027
rect 27077 25993 27111 26027
rect 27111 25993 27120 26027
rect 27068 25984 27120 25993
rect 27528 25984 27580 26036
rect 28448 25984 28500 26036
rect 8576 25916 8628 25968
rect 7840 25848 7892 25900
rect 23480 25848 23532 25900
rect 25504 25848 25556 25900
rect 26240 25848 26292 25900
rect 27988 25891 28040 25900
rect 27988 25857 27997 25891
rect 27997 25857 28031 25891
rect 28031 25857 28040 25891
rect 27988 25848 28040 25857
rect 28172 25891 28224 25900
rect 28172 25857 28181 25891
rect 28181 25857 28215 25891
rect 28215 25857 28224 25891
rect 28172 25848 28224 25857
rect 28356 25848 28408 25900
rect 29000 25848 29052 25900
rect 8576 25823 8628 25832
rect 8576 25789 8585 25823
rect 8585 25789 8619 25823
rect 8619 25789 8628 25823
rect 8576 25780 8628 25789
rect 9496 25823 9548 25832
rect 9496 25789 9505 25823
rect 9505 25789 9539 25823
rect 9539 25789 9548 25823
rect 9496 25780 9548 25789
rect 23204 25780 23256 25832
rect 24860 25823 24912 25832
rect 24860 25789 24869 25823
rect 24869 25789 24903 25823
rect 24903 25789 24912 25823
rect 24860 25780 24912 25789
rect 28908 25780 28960 25832
rect 29092 25823 29144 25832
rect 29092 25789 29101 25823
rect 29101 25789 29135 25823
rect 29135 25789 29144 25823
rect 29092 25780 29144 25789
rect 3056 25712 3108 25764
rect 28724 25712 28776 25764
rect 30564 25891 30616 25900
rect 30564 25857 30573 25891
rect 30573 25857 30607 25891
rect 30607 25857 30616 25891
rect 30564 25848 30616 25857
rect 34428 25984 34480 26036
rect 39856 25984 39908 26036
rect 33416 25959 33468 25968
rect 33416 25925 33425 25959
rect 33425 25925 33459 25959
rect 33459 25925 33468 25959
rect 33416 25916 33468 25925
rect 31116 25891 31168 25900
rect 31116 25857 31125 25891
rect 31125 25857 31159 25891
rect 31159 25857 31168 25891
rect 31116 25848 31168 25857
rect 29920 25780 29972 25832
rect 32404 25780 32456 25832
rect 33140 25848 33192 25900
rect 33600 25780 33652 25832
rect 32680 25755 32732 25764
rect 22468 25687 22520 25696
rect 22468 25653 22477 25687
rect 22477 25653 22511 25687
rect 22511 25653 22520 25687
rect 22468 25644 22520 25653
rect 28908 25644 28960 25696
rect 29460 25644 29512 25696
rect 31300 25687 31352 25696
rect 31300 25653 31309 25687
rect 31309 25653 31343 25687
rect 31343 25653 31352 25687
rect 31300 25644 31352 25653
rect 32680 25721 32689 25755
rect 32689 25721 32723 25755
rect 32723 25721 32732 25755
rect 32680 25712 32732 25721
rect 41880 25916 41932 25968
rect 44272 25916 44324 25968
rect 36452 25891 36504 25900
rect 36452 25857 36461 25891
rect 36461 25857 36495 25891
rect 36495 25857 36504 25891
rect 36452 25848 36504 25857
rect 39028 25891 39080 25900
rect 39028 25857 39037 25891
rect 39037 25857 39071 25891
rect 39071 25857 39080 25891
rect 39028 25848 39080 25857
rect 41604 25848 41656 25900
rect 44732 25780 44784 25832
rect 45008 25848 45060 25900
rect 45284 25848 45336 25900
rect 45744 25848 45796 25900
rect 46940 25848 46992 25900
rect 33600 25687 33652 25696
rect 33600 25653 33609 25687
rect 33609 25653 33643 25687
rect 33643 25653 33652 25687
rect 33600 25644 33652 25653
rect 33876 25644 33928 25696
rect 36544 25687 36596 25696
rect 36544 25653 36553 25687
rect 36553 25653 36587 25687
rect 36587 25653 36596 25687
rect 36544 25644 36596 25653
rect 38936 25644 38988 25696
rect 39948 25644 40000 25696
rect 44364 25644 44416 25696
rect 45376 25644 45428 25696
rect 45468 25644 45520 25696
rect 46480 25644 46532 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 25504 25483 25556 25492
rect 25504 25449 25513 25483
rect 25513 25449 25547 25483
rect 25547 25449 25556 25483
rect 25504 25440 25556 25449
rect 2136 25279 2188 25288
rect 2136 25245 2145 25279
rect 2145 25245 2179 25279
rect 2179 25245 2188 25279
rect 2136 25236 2188 25245
rect 18788 25304 18840 25356
rect 7840 25279 7892 25288
rect 7840 25245 7849 25279
rect 7849 25245 7883 25279
rect 7883 25245 7892 25279
rect 7840 25236 7892 25245
rect 12532 25236 12584 25288
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 22652 25279 22704 25288
rect 22652 25245 22661 25279
rect 22661 25245 22695 25279
rect 22695 25245 22704 25279
rect 22652 25236 22704 25245
rect 23112 25236 23164 25288
rect 23480 25279 23532 25288
rect 23480 25245 23489 25279
rect 23489 25245 23523 25279
rect 23523 25245 23532 25279
rect 23480 25236 23532 25245
rect 25136 25279 25188 25288
rect 25136 25245 25145 25279
rect 25145 25245 25179 25279
rect 25179 25245 25188 25279
rect 25136 25236 25188 25245
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 27620 25304 27672 25356
rect 26240 25279 26292 25288
rect 26240 25245 26249 25279
rect 26249 25245 26283 25279
rect 26283 25245 26292 25279
rect 26240 25236 26292 25245
rect 29092 25440 29144 25492
rect 31116 25440 31168 25492
rect 33324 25440 33376 25492
rect 36544 25440 36596 25492
rect 40316 25440 40368 25492
rect 44364 25483 44416 25492
rect 28724 25372 28776 25424
rect 29644 25415 29696 25424
rect 29644 25381 29653 25415
rect 29653 25381 29687 25415
rect 29687 25381 29696 25415
rect 29644 25372 29696 25381
rect 30380 25372 30432 25424
rect 35808 25415 35860 25424
rect 35808 25381 35817 25415
rect 35817 25381 35851 25415
rect 35851 25381 35860 25415
rect 35808 25372 35860 25381
rect 44364 25449 44373 25483
rect 44373 25449 44407 25483
rect 44407 25449 44416 25483
rect 44364 25440 44416 25449
rect 28540 25236 28592 25288
rect 28724 25279 28776 25288
rect 28724 25245 28733 25279
rect 28733 25245 28767 25279
rect 28767 25245 28776 25279
rect 28724 25236 28776 25245
rect 28908 25279 28960 25288
rect 28908 25245 28917 25279
rect 28917 25245 28951 25279
rect 28951 25245 28960 25279
rect 28908 25236 28960 25245
rect 41604 25304 41656 25356
rect 29460 25236 29512 25288
rect 32312 25236 32364 25288
rect 35900 25236 35952 25288
rect 35992 25279 36044 25288
rect 35992 25245 36001 25279
rect 36001 25245 36035 25279
rect 36035 25245 36044 25279
rect 40960 25279 41012 25288
rect 35992 25236 36044 25245
rect 40960 25245 40969 25279
rect 40969 25245 41003 25279
rect 41003 25245 41012 25279
rect 40960 25236 41012 25245
rect 44272 25304 44324 25356
rect 44180 25279 44232 25288
rect 44180 25245 44189 25279
rect 44189 25245 44223 25279
rect 44223 25245 44232 25279
rect 45284 25372 45336 25424
rect 45468 25372 45520 25424
rect 44548 25304 44600 25356
rect 44180 25236 44232 25245
rect 45376 25279 45428 25288
rect 29736 25168 29788 25220
rect 31300 25168 31352 25220
rect 36452 25168 36504 25220
rect 43444 25168 43496 25220
rect 45376 25245 45385 25279
rect 45385 25245 45419 25279
rect 45419 25245 45428 25279
rect 45376 25236 45428 25245
rect 46480 25347 46532 25356
rect 46480 25313 46489 25347
rect 46489 25313 46523 25347
rect 46523 25313 46532 25347
rect 46480 25304 46532 25313
rect 46756 25347 46808 25356
rect 46756 25313 46765 25347
rect 46765 25313 46799 25347
rect 46799 25313 46808 25347
rect 46756 25304 46808 25313
rect 45560 25168 45612 25220
rect 47768 25168 47820 25220
rect 2320 25100 2372 25152
rect 22744 25100 22796 25152
rect 22928 25100 22980 25152
rect 23296 25100 23348 25152
rect 27804 25100 27856 25152
rect 28632 25100 28684 25152
rect 41420 25100 41472 25152
rect 44916 25100 44968 25152
rect 45192 25100 45244 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 28724 24896 28776 24948
rect 33692 24896 33744 24948
rect 40960 24896 41012 24948
rect 2320 24871 2372 24880
rect 2320 24837 2329 24871
rect 2329 24837 2363 24871
rect 2363 24837 2372 24871
rect 2320 24828 2372 24837
rect 27620 24828 27672 24880
rect 2136 24803 2188 24812
rect 2136 24769 2145 24803
rect 2145 24769 2179 24803
rect 2179 24769 2188 24803
rect 2136 24760 2188 24769
rect 7840 24803 7892 24812
rect 7840 24769 7849 24803
rect 7849 24769 7883 24803
rect 7883 24769 7892 24803
rect 7840 24760 7892 24769
rect 23480 24760 23532 24812
rect 24768 24803 24820 24812
rect 24768 24769 24777 24803
rect 24777 24769 24811 24803
rect 24811 24769 24820 24803
rect 24768 24760 24820 24769
rect 27804 24803 27856 24812
rect 27804 24769 27813 24803
rect 27813 24769 27847 24803
rect 27847 24769 27856 24803
rect 27804 24760 27856 24769
rect 28632 24803 28684 24812
rect 28632 24769 28641 24803
rect 28641 24769 28675 24803
rect 28675 24769 28684 24803
rect 28632 24760 28684 24769
rect 32220 24760 32272 24812
rect 35716 24760 35768 24812
rect 37280 24760 37332 24812
rect 38752 24828 38804 24880
rect 39488 24760 39540 24812
rect 39580 24760 39632 24812
rect 2780 24735 2832 24744
rect 2780 24701 2789 24735
rect 2789 24701 2823 24735
rect 2823 24701 2832 24735
rect 2780 24692 2832 24701
rect 8024 24735 8076 24744
rect 8024 24701 8033 24735
rect 8033 24701 8067 24735
rect 8067 24701 8076 24735
rect 8024 24692 8076 24701
rect 22008 24735 22060 24744
rect 22008 24701 22017 24735
rect 22017 24701 22051 24735
rect 22051 24701 22060 24735
rect 22008 24692 22060 24701
rect 22192 24735 22244 24744
rect 22192 24701 22201 24735
rect 22201 24701 22235 24735
rect 22235 24701 22244 24735
rect 22192 24692 22244 24701
rect 3424 24624 3476 24676
rect 28356 24692 28408 24744
rect 29920 24692 29972 24744
rect 33416 24692 33468 24744
rect 33968 24692 34020 24744
rect 35532 24692 35584 24744
rect 35900 24624 35952 24676
rect 39120 24692 39172 24744
rect 43260 24760 43312 24812
rect 44180 24803 44232 24812
rect 44180 24769 44189 24803
rect 44189 24769 44223 24803
rect 44223 24769 44232 24803
rect 44180 24760 44232 24769
rect 44364 24828 44416 24880
rect 45560 24828 45612 24880
rect 44548 24803 44600 24812
rect 44548 24769 44557 24803
rect 44557 24769 44591 24803
rect 44591 24769 44600 24803
rect 44548 24760 44600 24769
rect 45284 24760 45336 24812
rect 45468 24803 45520 24812
rect 45468 24769 45477 24803
rect 45477 24769 45511 24803
rect 45511 24769 45520 24803
rect 45468 24760 45520 24769
rect 47032 24760 47084 24812
rect 47768 24803 47820 24812
rect 47768 24769 47777 24803
rect 47777 24769 47811 24803
rect 47811 24769 47820 24803
rect 47768 24760 47820 24769
rect 44364 24735 44416 24744
rect 44364 24701 44373 24735
rect 44373 24701 44407 24735
rect 44407 24701 44416 24735
rect 44364 24692 44416 24701
rect 38016 24624 38068 24676
rect 24952 24556 25004 24608
rect 31852 24556 31904 24608
rect 34796 24556 34848 24608
rect 37188 24556 37240 24608
rect 45560 24624 45612 24676
rect 39396 24599 39448 24608
rect 39396 24565 39405 24599
rect 39405 24565 39439 24599
rect 39439 24565 39448 24599
rect 39396 24556 39448 24565
rect 40592 24556 40644 24608
rect 44732 24599 44784 24608
rect 44732 24565 44741 24599
rect 44741 24565 44775 24599
rect 44775 24565 44784 24599
rect 44732 24556 44784 24565
rect 45468 24556 45520 24608
rect 45836 24556 45888 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 22192 24352 22244 24404
rect 23296 24395 23348 24404
rect 23296 24361 23305 24395
rect 23305 24361 23339 24395
rect 23339 24361 23348 24395
rect 23296 24352 23348 24361
rect 21916 24216 21968 24268
rect 33692 24352 33744 24404
rect 39120 24352 39172 24404
rect 39488 24352 39540 24404
rect 2044 24148 2096 24200
rect 22928 24191 22980 24200
rect 22928 24157 22937 24191
rect 22937 24157 22971 24191
rect 22971 24157 22980 24191
rect 22928 24148 22980 24157
rect 23940 24148 23992 24200
rect 28816 24148 28868 24200
rect 32128 24284 32180 24336
rect 33140 24284 33192 24336
rect 33968 24284 34020 24336
rect 31116 24216 31168 24268
rect 31484 24191 31536 24200
rect 31484 24157 31493 24191
rect 31493 24157 31527 24191
rect 31527 24157 31536 24191
rect 31484 24148 31536 24157
rect 32312 24216 32364 24268
rect 34520 24216 34572 24268
rect 35440 24216 35492 24268
rect 38016 24216 38068 24268
rect 40040 24284 40092 24336
rect 31668 24148 31720 24200
rect 31852 24191 31904 24200
rect 31852 24157 31861 24191
rect 31861 24157 31895 24191
rect 31895 24157 31904 24191
rect 31852 24148 31904 24157
rect 33140 24191 33192 24200
rect 22744 24080 22796 24132
rect 23112 24055 23164 24064
rect 23112 24021 23121 24055
rect 23121 24021 23155 24055
rect 23155 24021 23164 24055
rect 23112 24012 23164 24021
rect 24860 24080 24912 24132
rect 27804 24123 27856 24132
rect 27804 24089 27813 24123
rect 27813 24089 27847 24123
rect 27847 24089 27856 24123
rect 27804 24080 27856 24089
rect 28724 24080 28776 24132
rect 24768 24012 24820 24064
rect 27988 24055 28040 24064
rect 27988 24021 27997 24055
rect 27997 24021 28031 24055
rect 28031 24021 28040 24055
rect 27988 24012 28040 24021
rect 30840 24012 30892 24064
rect 32772 24055 32824 24064
rect 32772 24021 32781 24055
rect 32781 24021 32815 24055
rect 32815 24021 32824 24055
rect 32772 24012 32824 24021
rect 33140 24157 33149 24191
rect 33149 24157 33183 24191
rect 33183 24157 33192 24191
rect 33140 24148 33192 24157
rect 33600 24148 33652 24200
rect 33968 24191 34020 24200
rect 33968 24157 33977 24191
rect 33977 24157 34011 24191
rect 34011 24157 34020 24191
rect 33968 24148 34020 24157
rect 34796 24148 34848 24200
rect 35808 24191 35860 24200
rect 35808 24157 35842 24191
rect 35842 24157 35860 24191
rect 33324 24080 33376 24132
rect 35808 24148 35860 24157
rect 38660 24216 38712 24268
rect 39396 24216 39448 24268
rect 41420 24259 41472 24268
rect 41420 24225 41429 24259
rect 41429 24225 41463 24259
rect 41463 24225 41472 24259
rect 46204 24284 46256 24336
rect 41420 24216 41472 24225
rect 43904 24216 43956 24268
rect 38476 24148 38528 24200
rect 36268 24080 36320 24132
rect 38200 24123 38252 24132
rect 38200 24089 38209 24123
rect 38209 24089 38243 24123
rect 38243 24089 38252 24123
rect 38200 24080 38252 24089
rect 38384 24080 38436 24132
rect 39764 24148 39816 24200
rect 41236 24191 41288 24200
rect 34796 24012 34848 24064
rect 35348 24012 35400 24064
rect 36176 24012 36228 24064
rect 37280 24012 37332 24064
rect 37740 24012 37792 24064
rect 38844 24012 38896 24064
rect 41236 24157 41245 24191
rect 41245 24157 41279 24191
rect 41279 24157 41288 24191
rect 41236 24148 41288 24157
rect 43996 24191 44048 24200
rect 43996 24157 44005 24191
rect 44005 24157 44039 24191
rect 44039 24157 44048 24191
rect 43996 24148 44048 24157
rect 44732 24080 44784 24132
rect 47768 24216 47820 24268
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 45468 24191 45520 24200
rect 45468 24157 45477 24191
rect 45477 24157 45511 24191
rect 45511 24157 45520 24191
rect 45468 24148 45520 24157
rect 46940 24080 46992 24132
rect 43812 24012 43864 24064
rect 45100 24012 45152 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 22008 23808 22060 23860
rect 2044 23715 2096 23724
rect 2044 23681 2053 23715
rect 2053 23681 2087 23715
rect 2087 23681 2096 23715
rect 2044 23672 2096 23681
rect 2228 23647 2280 23656
rect 2228 23613 2237 23647
rect 2237 23613 2271 23647
rect 2271 23613 2280 23647
rect 2228 23604 2280 23613
rect 2780 23647 2832 23656
rect 2780 23613 2789 23647
rect 2789 23613 2823 23647
rect 2823 23613 2832 23647
rect 2780 23604 2832 23613
rect 23940 23647 23992 23656
rect 23940 23613 23949 23647
rect 23949 23613 23983 23647
rect 23983 23613 23992 23647
rect 23940 23604 23992 23613
rect 24308 23647 24360 23656
rect 24308 23613 24317 23647
rect 24317 23613 24351 23647
rect 24351 23613 24360 23647
rect 24308 23604 24360 23613
rect 24952 23672 25004 23724
rect 24584 23604 24636 23656
rect 27528 23808 27580 23860
rect 30380 23808 30432 23860
rect 31208 23740 31260 23792
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 25780 23715 25832 23724
rect 25780 23681 25786 23715
rect 25786 23681 25820 23715
rect 25820 23681 25832 23715
rect 25780 23672 25832 23681
rect 25964 23672 26016 23724
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 27160 23717 27212 23724
rect 27160 23683 27169 23717
rect 27169 23683 27203 23717
rect 27203 23683 27212 23717
rect 27160 23672 27212 23683
rect 27528 23715 27580 23724
rect 27528 23681 27537 23715
rect 27537 23681 27571 23715
rect 27571 23681 27580 23715
rect 30840 23715 30892 23724
rect 27528 23672 27580 23681
rect 30840 23681 30849 23715
rect 30849 23681 30883 23715
rect 30883 23681 30892 23715
rect 30840 23672 30892 23681
rect 31024 23715 31076 23724
rect 31024 23681 31033 23715
rect 31033 23681 31067 23715
rect 31067 23681 31076 23715
rect 31024 23672 31076 23681
rect 31116 23715 31168 23724
rect 31116 23681 31125 23715
rect 31125 23681 31159 23715
rect 31159 23681 31168 23715
rect 33600 23808 33652 23860
rect 35992 23808 36044 23860
rect 38384 23808 38436 23860
rect 38844 23851 38896 23860
rect 38844 23817 38853 23851
rect 38853 23817 38887 23851
rect 38887 23817 38896 23851
rect 38844 23808 38896 23817
rect 39580 23851 39632 23860
rect 39580 23817 39589 23851
rect 39589 23817 39623 23851
rect 39623 23817 39632 23851
rect 39580 23808 39632 23817
rect 43996 23808 44048 23860
rect 46940 23851 46992 23860
rect 46940 23817 46949 23851
rect 46949 23817 46983 23851
rect 46983 23817 46992 23851
rect 46940 23808 46992 23817
rect 32772 23783 32824 23792
rect 32772 23749 32806 23783
rect 32806 23749 32824 23783
rect 32772 23740 32824 23749
rect 36176 23783 36228 23792
rect 36176 23749 36185 23783
rect 36185 23749 36219 23783
rect 36219 23749 36228 23783
rect 36176 23740 36228 23749
rect 31116 23672 31168 23681
rect 32312 23672 32364 23724
rect 34428 23672 34480 23724
rect 34612 23715 34664 23724
rect 34612 23681 34646 23715
rect 34646 23681 34664 23715
rect 34612 23672 34664 23681
rect 35716 23672 35768 23724
rect 38568 23740 38620 23792
rect 26792 23536 26844 23588
rect 25688 23468 25740 23520
rect 26424 23468 26476 23520
rect 30748 23604 30800 23656
rect 38384 23536 38436 23588
rect 39856 23672 39908 23724
rect 42432 23740 42484 23792
rect 40592 23672 40644 23724
rect 43168 23672 43220 23724
rect 43260 23715 43312 23724
rect 43260 23681 43269 23715
rect 43269 23681 43303 23715
rect 43303 23681 43312 23715
rect 43904 23715 43956 23724
rect 43260 23672 43312 23681
rect 40040 23604 40092 23656
rect 42800 23604 42852 23656
rect 43904 23681 43913 23715
rect 43913 23681 43947 23715
rect 43947 23681 43956 23715
rect 43904 23672 43956 23681
rect 45836 23672 45888 23724
rect 46020 23715 46072 23724
rect 46020 23681 46029 23715
rect 46029 23681 46063 23715
rect 46063 23681 46072 23715
rect 46020 23672 46072 23681
rect 46112 23715 46164 23724
rect 46112 23681 46121 23715
rect 46121 23681 46155 23715
rect 46155 23681 46164 23715
rect 46112 23672 46164 23681
rect 46296 23715 46348 23724
rect 46296 23681 46305 23715
rect 46305 23681 46339 23715
rect 46339 23681 46348 23715
rect 46296 23672 46348 23681
rect 47216 23672 47268 23724
rect 47768 23715 47820 23724
rect 47768 23681 47777 23715
rect 47777 23681 47811 23715
rect 47811 23681 47820 23715
rect 47768 23672 47820 23681
rect 43812 23647 43864 23656
rect 43812 23613 43821 23647
rect 43821 23613 43855 23647
rect 43855 23613 43864 23647
rect 43812 23604 43864 23613
rect 29552 23468 29604 23520
rect 30012 23468 30064 23520
rect 35532 23468 35584 23520
rect 36636 23468 36688 23520
rect 38476 23468 38528 23520
rect 45008 23536 45060 23588
rect 39856 23468 39908 23520
rect 46940 23468 46992 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2228 23264 2280 23316
rect 24308 23264 24360 23316
rect 26976 23264 27028 23316
rect 32312 23264 32364 23316
rect 34612 23264 34664 23316
rect 35716 23264 35768 23316
rect 24584 23196 24636 23248
rect 22100 23128 22152 23180
rect 2228 23060 2280 23112
rect 16948 23060 17000 23112
rect 25780 23128 25832 23180
rect 24952 23103 25004 23112
rect 24952 23069 24961 23103
rect 24961 23069 24995 23103
rect 24995 23069 25004 23103
rect 24952 23060 25004 23069
rect 30472 23239 30524 23248
rect 30472 23205 30481 23239
rect 30481 23205 30515 23239
rect 30515 23205 30524 23239
rect 30472 23196 30524 23205
rect 30656 23196 30708 23248
rect 36912 23264 36964 23316
rect 41144 23264 41196 23316
rect 41236 23264 41288 23316
rect 46112 23264 46164 23316
rect 47032 23264 47084 23316
rect 39764 23196 39816 23248
rect 27988 23128 28040 23180
rect 30012 23128 30064 23180
rect 28724 23103 28776 23112
rect 25780 22992 25832 23044
rect 26792 22992 26844 23044
rect 27160 22924 27212 22976
rect 27436 22924 27488 22976
rect 28724 23069 28733 23103
rect 28733 23069 28767 23103
rect 28767 23069 28776 23103
rect 28724 23060 28776 23069
rect 28816 23103 28868 23112
rect 28816 23069 28830 23103
rect 28830 23069 28864 23103
rect 28864 23069 28868 23103
rect 28816 23060 28868 23069
rect 30564 23060 30616 23112
rect 31024 23060 31076 23112
rect 31208 23103 31260 23112
rect 31208 23069 31217 23103
rect 31217 23069 31251 23103
rect 31251 23069 31260 23103
rect 39028 23128 39080 23180
rect 31208 23060 31260 23069
rect 35348 23060 35400 23112
rect 35532 23103 35584 23112
rect 35532 23069 35541 23103
rect 35541 23069 35575 23103
rect 35575 23069 35584 23103
rect 35532 23060 35584 23069
rect 36452 23060 36504 23112
rect 37740 23103 37792 23112
rect 37740 23069 37749 23103
rect 37749 23069 37783 23103
rect 37783 23069 37792 23103
rect 37740 23060 37792 23069
rect 39856 23103 39908 23112
rect 39856 23069 39865 23103
rect 39865 23069 39899 23103
rect 39899 23069 39908 23103
rect 39856 23060 39908 23069
rect 39948 23060 40000 23112
rect 40592 23103 40644 23112
rect 40592 23069 40601 23103
rect 40601 23069 40635 23103
rect 40635 23069 40644 23103
rect 40592 23060 40644 23069
rect 40776 23103 40828 23112
rect 40776 23069 40785 23103
rect 40785 23069 40819 23103
rect 40819 23069 40828 23103
rect 40776 23060 40828 23069
rect 45008 23103 45060 23112
rect 30288 22992 30340 23044
rect 30380 22924 30432 22976
rect 30564 22924 30616 22976
rect 40040 22992 40092 23044
rect 35900 22924 35952 22976
rect 39488 22924 39540 22976
rect 39580 22924 39632 22976
rect 40132 22924 40184 22976
rect 45008 23069 45017 23103
rect 45017 23069 45051 23103
rect 45051 23069 45060 23103
rect 45008 23060 45060 23069
rect 45284 23060 45336 23112
rect 45652 23060 45704 23112
rect 46664 23103 46716 23112
rect 46664 23069 46673 23103
rect 46673 23069 46707 23103
rect 46707 23069 46716 23103
rect 46664 23060 46716 23069
rect 46940 23103 46992 23112
rect 46940 23069 46974 23103
rect 46974 23069 46992 23103
rect 46940 23060 46992 23069
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 17868 22720 17920 22772
rect 30656 22720 30708 22772
rect 31024 22720 31076 22772
rect 31484 22720 31536 22772
rect 23940 22652 23992 22704
rect 30288 22652 30340 22704
rect 24584 22627 24636 22636
rect 24584 22593 24593 22627
rect 24593 22593 24627 22627
rect 24627 22593 24636 22627
rect 24584 22584 24636 22593
rect 24676 22627 24728 22636
rect 24676 22593 24685 22627
rect 24685 22593 24719 22627
rect 24719 22593 24728 22627
rect 29552 22627 29604 22636
rect 24676 22584 24728 22593
rect 29552 22593 29561 22627
rect 29561 22593 29595 22627
rect 29595 22593 29604 22627
rect 29552 22584 29604 22593
rect 29828 22627 29880 22636
rect 29828 22593 29862 22627
rect 29862 22593 29880 22627
rect 29828 22584 29880 22593
rect 31668 22584 31720 22636
rect 33140 22720 33192 22772
rect 33416 22720 33468 22772
rect 35900 22695 35952 22704
rect 35900 22661 35909 22695
rect 35909 22661 35943 22695
rect 35943 22661 35952 22695
rect 35900 22652 35952 22661
rect 37188 22652 37240 22704
rect 39488 22695 39540 22704
rect 32588 22627 32640 22636
rect 32588 22593 32597 22627
rect 32597 22593 32631 22627
rect 32631 22593 32640 22627
rect 32588 22584 32640 22593
rect 35992 22584 36044 22636
rect 36544 22584 36596 22636
rect 36636 22584 36688 22636
rect 39488 22661 39497 22695
rect 39497 22661 39531 22695
rect 39531 22661 39540 22695
rect 39488 22652 39540 22661
rect 38660 22627 38712 22636
rect 38660 22593 38669 22627
rect 38669 22593 38703 22627
rect 38703 22593 38712 22627
rect 38660 22584 38712 22593
rect 40040 22720 40092 22772
rect 40776 22720 40828 22772
rect 41144 22720 41196 22772
rect 39948 22652 40000 22704
rect 32312 22516 32364 22568
rect 40132 22584 40184 22636
rect 40316 22627 40368 22636
rect 40316 22593 40325 22627
rect 40325 22593 40359 22627
rect 40359 22593 40368 22627
rect 40316 22584 40368 22593
rect 40408 22584 40460 22636
rect 45100 22652 45152 22704
rect 45376 22652 45428 22704
rect 39764 22516 39816 22568
rect 40592 22559 40644 22568
rect 40592 22525 40601 22559
rect 40601 22525 40635 22559
rect 40635 22525 40644 22559
rect 40592 22516 40644 22525
rect 42064 22584 42116 22636
rect 42432 22627 42484 22636
rect 42432 22593 42441 22627
rect 42441 22593 42475 22627
rect 42475 22593 42484 22627
rect 42432 22584 42484 22593
rect 42524 22584 42576 22636
rect 45008 22584 45060 22636
rect 24308 22380 24360 22432
rect 31208 22380 31260 22432
rect 36084 22380 36136 22432
rect 39120 22380 39172 22432
rect 41512 22448 41564 22500
rect 40408 22380 40460 22432
rect 44180 22380 44232 22432
rect 45652 22423 45704 22432
rect 45652 22389 45661 22423
rect 45661 22389 45695 22423
rect 45695 22389 45704 22423
rect 45652 22380 45704 22389
rect 47032 22423 47084 22432
rect 47032 22389 47041 22423
rect 47041 22389 47075 22423
rect 47075 22389 47084 22423
rect 47032 22380 47084 22389
rect 47676 22423 47728 22432
rect 47676 22389 47685 22423
rect 47685 22389 47719 22423
rect 47719 22389 47728 22423
rect 47676 22380 47728 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 25780 22219 25832 22228
rect 25780 22185 25789 22219
rect 25789 22185 25823 22219
rect 25823 22185 25832 22219
rect 25780 22176 25832 22185
rect 26424 22219 26476 22228
rect 26424 22185 26433 22219
rect 26433 22185 26467 22219
rect 26467 22185 26476 22219
rect 26424 22176 26476 22185
rect 26976 22176 27028 22228
rect 29828 22176 29880 22228
rect 30380 22219 30432 22228
rect 30380 22185 30389 22219
rect 30389 22185 30423 22219
rect 30423 22185 30432 22219
rect 30380 22176 30432 22185
rect 31116 22176 31168 22228
rect 39120 22176 39172 22228
rect 39856 22176 39908 22228
rect 40316 22176 40368 22228
rect 42524 22176 42576 22228
rect 17224 22108 17276 22160
rect 17868 22108 17920 22160
rect 30472 22108 30524 22160
rect 27620 22040 27672 22092
rect 28356 22040 28408 22092
rect 29368 22040 29420 22092
rect 31024 22083 31076 22092
rect 2044 21972 2096 22024
rect 24768 21904 24820 21956
rect 24860 21904 24912 21956
rect 25780 21904 25832 21956
rect 27160 22015 27212 22024
rect 27160 21981 27169 22015
rect 27169 21981 27203 22015
rect 27203 21981 27212 22015
rect 31024 22049 31033 22083
rect 31033 22049 31067 22083
rect 31067 22049 31076 22083
rect 31024 22040 31076 22049
rect 31116 22040 31168 22092
rect 31760 22040 31812 22092
rect 32588 22083 32640 22092
rect 32588 22049 32597 22083
rect 32597 22049 32631 22083
rect 32631 22049 32640 22083
rect 32588 22040 32640 22049
rect 35440 22040 35492 22092
rect 27160 21972 27212 21981
rect 30564 21972 30616 22024
rect 31208 21972 31260 22024
rect 39580 21972 39632 22024
rect 26424 21879 26476 21888
rect 26424 21845 26449 21879
rect 26449 21845 26476 21879
rect 26608 21879 26660 21888
rect 26424 21836 26476 21845
rect 26608 21845 26617 21879
rect 26617 21845 26651 21879
rect 26651 21845 26660 21879
rect 26608 21836 26660 21845
rect 26700 21836 26752 21888
rect 34612 21904 34664 21956
rect 35900 21904 35952 21956
rect 41420 22040 41472 22092
rect 39948 22015 40000 22024
rect 39948 21981 39957 22015
rect 39957 21981 39991 22015
rect 39991 21981 40000 22015
rect 39948 21972 40000 21981
rect 40040 22015 40092 22024
rect 40040 21981 40050 22015
rect 40050 21981 40084 22015
rect 40084 21981 40092 22015
rect 40040 21972 40092 21981
rect 40408 22015 40460 22024
rect 40408 21981 40422 22015
rect 40422 21981 40456 22015
rect 40456 21981 40460 22015
rect 40408 21972 40460 21981
rect 40684 21972 40736 22024
rect 41788 21972 41840 22024
rect 39856 21904 39908 21956
rect 40592 21904 40644 21956
rect 41972 21981 41981 22002
rect 41981 21981 42015 22002
rect 42015 21981 42024 22002
rect 41972 21950 42024 21981
rect 42156 21972 42208 22024
rect 44180 22040 44232 22092
rect 45008 22040 45060 22092
rect 47032 22040 47084 22092
rect 48136 22083 48188 22092
rect 48136 22049 48145 22083
rect 48145 22049 48179 22083
rect 48179 22049 48188 22083
rect 48136 22040 48188 22049
rect 42984 21972 43036 22024
rect 42708 21904 42760 21956
rect 44548 21972 44600 22024
rect 45376 22015 45428 22024
rect 45376 21981 45385 22015
rect 45385 21981 45419 22015
rect 45419 21981 45428 22015
rect 45376 21972 45428 21981
rect 45468 22015 45520 22024
rect 45468 21981 45477 22015
rect 45477 21981 45511 22015
rect 45511 21981 45520 22015
rect 45468 21972 45520 21981
rect 44732 21904 44784 21956
rect 47676 21904 47728 21956
rect 27344 21879 27396 21888
rect 27344 21845 27353 21879
rect 27353 21845 27387 21879
rect 27387 21845 27396 21879
rect 27344 21836 27396 21845
rect 37188 21879 37240 21888
rect 37188 21845 37197 21879
rect 37197 21845 37231 21879
rect 37231 21845 37240 21879
rect 37188 21836 37240 21845
rect 39488 21836 39540 21888
rect 42616 21836 42668 21888
rect 42984 21879 43036 21888
rect 42984 21845 42993 21879
rect 42993 21845 43027 21879
rect 43027 21845 43036 21879
rect 42984 21836 43036 21845
rect 44272 21836 44324 21888
rect 45284 21836 45336 21888
rect 45560 21836 45612 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 24768 21632 24820 21684
rect 28816 21632 28868 21684
rect 30380 21675 30432 21684
rect 30380 21641 30405 21675
rect 30405 21641 30432 21675
rect 30380 21632 30432 21641
rect 35900 21675 35952 21684
rect 35900 21641 35909 21675
rect 35909 21641 35943 21675
rect 35943 21641 35952 21675
rect 35900 21632 35952 21641
rect 39948 21632 40000 21684
rect 41972 21632 42024 21684
rect 42984 21675 43036 21684
rect 42984 21641 42993 21675
rect 42993 21641 43027 21675
rect 43027 21641 43036 21675
rect 42984 21632 43036 21641
rect 44916 21632 44968 21684
rect 45284 21632 45336 21684
rect 2044 21539 2096 21548
rect 2044 21505 2053 21539
rect 2053 21505 2087 21539
rect 2087 21505 2096 21539
rect 2044 21496 2096 21505
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 24308 21496 24360 21505
rect 27344 21564 27396 21616
rect 2412 21428 2464 21480
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 2780 21428 2832 21437
rect 24584 21471 24636 21480
rect 24584 21437 24593 21471
rect 24593 21437 24627 21471
rect 24627 21437 24636 21471
rect 24584 21428 24636 21437
rect 2872 21360 2924 21412
rect 16764 21360 16816 21412
rect 24676 21360 24728 21412
rect 26608 21496 26660 21548
rect 30564 21564 30616 21616
rect 30656 21564 30708 21616
rect 31116 21564 31168 21616
rect 26424 21428 26476 21480
rect 28264 21496 28316 21548
rect 28448 21496 28500 21548
rect 31208 21539 31260 21548
rect 26976 21471 27028 21480
rect 26976 21437 26985 21471
rect 26985 21437 27019 21471
rect 27019 21437 27028 21471
rect 31208 21505 31217 21539
rect 31217 21505 31251 21539
rect 31251 21505 31260 21539
rect 31208 21496 31260 21505
rect 42708 21564 42760 21616
rect 34428 21539 34480 21548
rect 34428 21505 34437 21539
rect 34437 21505 34471 21539
rect 34471 21505 34480 21539
rect 34428 21496 34480 21505
rect 36084 21539 36136 21548
rect 36084 21505 36093 21539
rect 36093 21505 36127 21539
rect 36127 21505 36136 21539
rect 36084 21496 36136 21505
rect 36544 21496 36596 21548
rect 38108 21496 38160 21548
rect 38660 21539 38712 21548
rect 26976 21428 27028 21437
rect 24124 21335 24176 21344
rect 24124 21301 24133 21335
rect 24133 21301 24167 21335
rect 24167 21301 24176 21335
rect 24124 21292 24176 21301
rect 26240 21292 26292 21344
rect 27160 21292 27212 21344
rect 27988 21292 28040 21344
rect 37188 21428 37240 21480
rect 30288 21360 30340 21412
rect 33876 21360 33928 21412
rect 37924 21360 37976 21412
rect 38660 21505 38669 21539
rect 38669 21505 38703 21539
rect 38703 21505 38712 21539
rect 38660 21496 38712 21505
rect 38844 21539 38896 21548
rect 38844 21505 38853 21539
rect 38853 21505 38887 21539
rect 38887 21505 38896 21539
rect 38844 21496 38896 21505
rect 39488 21539 39540 21548
rect 39488 21505 39497 21539
rect 39497 21505 39531 21539
rect 39531 21505 39540 21539
rect 39488 21496 39540 21505
rect 39856 21539 39908 21548
rect 38568 21471 38620 21480
rect 38568 21437 38577 21471
rect 38577 21437 38611 21471
rect 38611 21437 38620 21471
rect 38568 21428 38620 21437
rect 39856 21505 39865 21539
rect 39865 21505 39899 21539
rect 39899 21505 39908 21539
rect 39856 21496 39908 21505
rect 40040 21539 40092 21548
rect 40040 21505 40049 21539
rect 40049 21505 40083 21539
rect 40083 21505 40092 21539
rect 40040 21496 40092 21505
rect 41880 21539 41932 21548
rect 39764 21471 39816 21480
rect 39764 21437 39773 21471
rect 39773 21437 39807 21471
rect 39807 21437 39816 21471
rect 41880 21505 41889 21539
rect 41889 21505 41923 21539
rect 41923 21505 41932 21539
rect 41880 21496 41932 21505
rect 44548 21564 44600 21616
rect 44732 21564 44784 21616
rect 42892 21496 42944 21548
rect 43076 21539 43128 21548
rect 43076 21505 43085 21539
rect 43085 21505 43119 21539
rect 43119 21505 43128 21539
rect 43076 21496 43128 21505
rect 44180 21539 44232 21548
rect 44180 21505 44189 21539
rect 44189 21505 44223 21539
rect 44223 21505 44232 21539
rect 44180 21496 44232 21505
rect 44916 21496 44968 21548
rect 45652 21496 45704 21548
rect 39764 21428 39816 21437
rect 44364 21428 44416 21480
rect 44548 21471 44600 21480
rect 44548 21437 44557 21471
rect 44557 21437 44591 21471
rect 44591 21437 44600 21471
rect 44548 21428 44600 21437
rect 45100 21428 45152 21480
rect 48136 21496 48188 21548
rect 47676 21471 47728 21480
rect 47676 21437 47685 21471
rect 47685 21437 47719 21471
rect 47719 21437 47728 21471
rect 47676 21428 47728 21437
rect 28632 21335 28684 21344
rect 28632 21301 28641 21335
rect 28641 21301 28675 21335
rect 28675 21301 28684 21335
rect 28632 21292 28684 21301
rect 30656 21292 30708 21344
rect 31024 21335 31076 21344
rect 31024 21301 31033 21335
rect 31033 21301 31067 21335
rect 31067 21301 31076 21335
rect 31024 21292 31076 21301
rect 38568 21292 38620 21344
rect 43260 21292 43312 21344
rect 45008 21292 45060 21344
rect 46112 21292 46164 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2412 21131 2464 21140
rect 2412 21097 2421 21131
rect 2421 21097 2455 21131
rect 2455 21097 2464 21131
rect 2412 21088 2464 21097
rect 24584 21088 24636 21140
rect 27988 21088 28040 21140
rect 28816 21088 28868 21140
rect 31576 21088 31628 21140
rect 38108 21131 38160 21140
rect 38108 21097 38117 21131
rect 38117 21097 38151 21131
rect 38151 21097 38160 21131
rect 38108 21088 38160 21097
rect 39764 21088 39816 21140
rect 43076 21088 43128 21140
rect 45100 21131 45152 21140
rect 45100 21097 45109 21131
rect 45109 21097 45143 21131
rect 45143 21097 45152 21131
rect 45100 21088 45152 21097
rect 45192 21088 45244 21140
rect 47676 21088 47728 21140
rect 48136 21131 48188 21140
rect 48136 21097 48145 21131
rect 48145 21097 48179 21131
rect 48179 21097 48188 21131
rect 48136 21088 48188 21097
rect 27620 21020 27672 21072
rect 33324 21020 33376 21072
rect 39120 21020 39172 21072
rect 41788 21020 41840 21072
rect 44364 21020 44416 21072
rect 44824 21020 44876 21072
rect 29552 20952 29604 21004
rect 29920 20995 29972 21004
rect 29920 20961 29929 20995
rect 29929 20961 29963 20995
rect 29963 20961 29972 20995
rect 29920 20952 29972 20961
rect 31208 20952 31260 21004
rect 2872 20884 2924 20936
rect 3148 20927 3200 20936
rect 3148 20893 3157 20927
rect 3157 20893 3191 20927
rect 3191 20893 3200 20927
rect 3148 20884 3200 20893
rect 26240 20927 26292 20936
rect 26240 20893 26249 20927
rect 26249 20893 26283 20927
rect 26283 20893 26292 20927
rect 26240 20884 26292 20893
rect 26700 20884 26752 20936
rect 27344 20884 27396 20936
rect 31760 20927 31812 20936
rect 24124 20816 24176 20868
rect 24860 20816 24912 20868
rect 31760 20893 31769 20927
rect 31769 20893 31803 20927
rect 31803 20893 31812 20927
rect 31760 20884 31812 20893
rect 34612 20952 34664 21004
rect 33876 20927 33928 20936
rect 33876 20893 33885 20927
rect 33885 20893 33919 20927
rect 33919 20893 33928 20927
rect 33876 20884 33928 20893
rect 34796 20884 34848 20936
rect 34980 20884 35032 20936
rect 35624 20927 35676 20936
rect 35624 20893 35633 20927
rect 35633 20893 35667 20927
rect 35667 20893 35676 20927
rect 35624 20884 35676 20893
rect 37464 20927 37516 20936
rect 37464 20893 37473 20927
rect 37473 20893 37507 20927
rect 37507 20893 37516 20927
rect 37464 20884 37516 20893
rect 38200 20952 38252 21004
rect 38844 20952 38896 21004
rect 37924 20927 37976 20936
rect 37924 20893 37938 20927
rect 37938 20893 37972 20927
rect 37972 20893 37976 20927
rect 39028 20927 39080 20936
rect 37924 20884 37976 20893
rect 39028 20893 39037 20927
rect 39037 20893 39071 20927
rect 39071 20893 39080 20927
rect 39028 20884 39080 20893
rect 39304 20927 39356 20936
rect 39304 20893 39313 20927
rect 39313 20893 39347 20927
rect 39347 20893 39356 20927
rect 39304 20884 39356 20893
rect 39580 20952 39632 21004
rect 44732 20952 44784 21004
rect 46756 20995 46808 21004
rect 42984 20884 43036 20936
rect 45008 20927 45060 20936
rect 45008 20893 45017 20927
rect 45017 20893 45051 20927
rect 45051 20893 45060 20927
rect 45008 20884 45060 20893
rect 45376 20884 45428 20936
rect 46756 20961 46765 20995
rect 46765 20961 46799 20995
rect 46799 20961 46808 20995
rect 46756 20952 46808 20961
rect 46020 20927 46072 20936
rect 46020 20893 46029 20927
rect 46029 20893 46063 20927
rect 46063 20893 46072 20927
rect 46020 20884 46072 20893
rect 46112 20927 46164 20936
rect 46112 20893 46121 20927
rect 46121 20893 46155 20927
rect 46155 20893 46164 20927
rect 46112 20884 46164 20893
rect 46296 20927 46348 20936
rect 46296 20893 46305 20927
rect 46305 20893 46339 20927
rect 46339 20893 46348 20927
rect 46296 20884 46348 20893
rect 28632 20816 28684 20868
rect 37740 20859 37792 20868
rect 37740 20825 37749 20859
rect 37749 20825 37783 20859
rect 37783 20825 37792 20859
rect 37740 20816 37792 20825
rect 38568 20816 38620 20868
rect 26240 20748 26292 20800
rect 27068 20748 27120 20800
rect 34428 20748 34480 20800
rect 38660 20748 38712 20800
rect 41420 20816 41472 20868
rect 39488 20748 39540 20800
rect 42708 20748 42760 20800
rect 42892 20748 42944 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 28448 20587 28500 20596
rect 28448 20553 28457 20587
rect 28457 20553 28491 20587
rect 28491 20553 28500 20587
rect 28448 20544 28500 20553
rect 30656 20544 30708 20596
rect 3148 20476 3200 20528
rect 27344 20519 27396 20528
rect 27344 20485 27353 20519
rect 27353 20485 27387 20519
rect 27387 20485 27396 20519
rect 27344 20476 27396 20485
rect 28264 20476 28316 20528
rect 34704 20544 34756 20596
rect 34796 20544 34848 20596
rect 26240 20408 26292 20460
rect 26332 20451 26384 20460
rect 26332 20417 26341 20451
rect 26341 20417 26375 20451
rect 26375 20417 26384 20451
rect 26332 20408 26384 20417
rect 26976 20408 27028 20460
rect 2596 20340 2648 20392
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 26424 20272 26476 20324
rect 27252 20272 27304 20324
rect 28816 20408 28868 20460
rect 29920 20451 29972 20460
rect 29920 20417 29929 20451
rect 29929 20417 29963 20451
rect 29963 20417 29972 20451
rect 29920 20408 29972 20417
rect 30196 20451 30248 20460
rect 30196 20417 30230 20451
rect 30230 20417 30248 20451
rect 33232 20451 33284 20460
rect 30196 20408 30248 20417
rect 33232 20417 33241 20451
rect 33241 20417 33275 20451
rect 33275 20417 33284 20451
rect 33232 20408 33284 20417
rect 33416 20408 33468 20460
rect 35440 20476 35492 20528
rect 37464 20544 37516 20596
rect 37740 20544 37792 20596
rect 39304 20544 39356 20596
rect 41696 20544 41748 20596
rect 41880 20544 41932 20596
rect 45468 20544 45520 20596
rect 28356 20340 28408 20392
rect 31760 20340 31812 20392
rect 33876 20408 33928 20460
rect 34980 20408 35032 20460
rect 37464 20408 37516 20460
rect 42156 20476 42208 20528
rect 45560 20476 45612 20528
rect 37188 20340 37240 20392
rect 37832 20408 37884 20460
rect 39120 20451 39172 20460
rect 39120 20417 39129 20451
rect 39129 20417 39163 20451
rect 39163 20417 39172 20451
rect 39120 20408 39172 20417
rect 38200 20340 38252 20392
rect 39488 20408 39540 20460
rect 44824 20451 44876 20460
rect 44824 20417 44833 20451
rect 44833 20417 44867 20451
rect 44867 20417 44876 20451
rect 44824 20408 44876 20417
rect 44916 20408 44968 20460
rect 46572 20408 46624 20460
rect 44732 20340 44784 20392
rect 25872 20247 25924 20256
rect 25872 20213 25881 20247
rect 25881 20213 25915 20247
rect 25915 20213 25924 20247
rect 25872 20204 25924 20213
rect 35348 20272 35400 20324
rect 38384 20272 38436 20324
rect 28264 20247 28316 20256
rect 28264 20213 28273 20247
rect 28273 20213 28307 20247
rect 28307 20213 28316 20247
rect 28264 20204 28316 20213
rect 30288 20204 30340 20256
rect 33692 20204 33744 20256
rect 34704 20204 34756 20256
rect 35624 20204 35676 20256
rect 36360 20204 36412 20256
rect 41880 20204 41932 20256
rect 46480 20204 46532 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2596 20043 2648 20052
rect 2596 20009 2605 20043
rect 2605 20009 2639 20043
rect 2639 20009 2648 20043
rect 2596 20000 2648 20009
rect 26332 20000 26384 20052
rect 27344 20000 27396 20052
rect 30196 20043 30248 20052
rect 30196 20009 30205 20043
rect 30205 20009 30239 20043
rect 30239 20009 30248 20043
rect 30196 20000 30248 20009
rect 33876 20000 33928 20052
rect 31024 19932 31076 19984
rect 33692 19975 33744 19984
rect 33692 19941 33701 19975
rect 33701 19941 33735 19975
rect 33735 19941 33744 19975
rect 33692 19932 33744 19941
rect 24860 19907 24912 19916
rect 24860 19873 24869 19907
rect 24869 19873 24903 19907
rect 24903 19873 24912 19907
rect 24860 19864 24912 19873
rect 31760 19907 31812 19916
rect 31760 19873 31769 19907
rect 31769 19873 31803 19907
rect 31803 19873 31812 19907
rect 31760 19864 31812 19873
rect 33232 19864 33284 19916
rect 34428 19864 34480 19916
rect 17316 19796 17368 19848
rect 30288 19796 30340 19848
rect 31852 19796 31904 19848
rect 32496 19796 32548 19848
rect 35348 20000 35400 20052
rect 37464 20043 37516 20052
rect 37464 20009 37473 20043
rect 37473 20009 37507 20043
rect 37507 20009 37516 20043
rect 37464 20000 37516 20009
rect 40500 20000 40552 20052
rect 41512 20000 41564 20052
rect 45468 20000 45520 20052
rect 35440 19864 35492 19916
rect 36360 19839 36412 19848
rect 36360 19805 36394 19839
rect 36394 19805 36412 19839
rect 36360 19796 36412 19805
rect 38200 19975 38252 19984
rect 38200 19941 38209 19975
rect 38209 19941 38243 19975
rect 38243 19941 38252 19975
rect 38200 19932 38252 19941
rect 39304 19864 39356 19916
rect 42064 19907 42116 19916
rect 39120 19796 39172 19848
rect 39672 19796 39724 19848
rect 40224 19839 40276 19848
rect 40224 19805 40233 19839
rect 40233 19805 40267 19839
rect 40267 19805 40276 19839
rect 42064 19873 42073 19907
rect 42073 19873 42107 19907
rect 42107 19873 42116 19907
rect 42064 19864 42116 19873
rect 43260 19864 43312 19916
rect 44456 19864 44508 19916
rect 46480 19907 46532 19916
rect 46480 19873 46489 19907
rect 46489 19873 46523 19907
rect 46523 19873 46532 19907
rect 46480 19864 46532 19873
rect 48136 19907 48188 19916
rect 48136 19873 48145 19907
rect 48145 19873 48179 19907
rect 48179 19873 48188 19907
rect 48136 19864 48188 19873
rect 40224 19796 40276 19805
rect 44824 19796 44876 19848
rect 45284 19796 45336 19848
rect 25872 19728 25924 19780
rect 27160 19728 27212 19780
rect 32404 19728 32456 19780
rect 34704 19771 34756 19780
rect 34704 19737 34713 19771
rect 34713 19737 34747 19771
rect 34747 19737 34756 19771
rect 34704 19728 34756 19737
rect 37188 19728 37240 19780
rect 2504 19660 2556 19712
rect 32312 19660 32364 19712
rect 33416 19660 33468 19712
rect 34796 19660 34848 19712
rect 38844 19703 38896 19712
rect 38844 19669 38853 19703
rect 38853 19669 38887 19703
rect 38887 19669 38896 19703
rect 38844 19660 38896 19669
rect 40316 19728 40368 19780
rect 42340 19771 42392 19780
rect 42340 19737 42374 19771
rect 42374 19737 42392 19771
rect 42340 19728 42392 19737
rect 40868 19660 40920 19712
rect 45192 19728 45244 19780
rect 47768 19728 47820 19780
rect 42616 19660 42668 19712
rect 43628 19660 43680 19712
rect 44364 19703 44416 19712
rect 44364 19669 44373 19703
rect 44373 19669 44407 19703
rect 44407 19669 44416 19703
rect 44364 19660 44416 19669
rect 46296 19660 46348 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 27160 19499 27212 19508
rect 27160 19465 27169 19499
rect 27169 19465 27203 19499
rect 27203 19465 27212 19499
rect 27160 19456 27212 19465
rect 32404 19499 32456 19508
rect 32404 19465 32413 19499
rect 32413 19465 32447 19499
rect 32447 19465 32456 19499
rect 32404 19456 32456 19465
rect 34428 19499 34480 19508
rect 34428 19465 34437 19499
rect 34437 19465 34471 19499
rect 34471 19465 34480 19499
rect 34428 19456 34480 19465
rect 37832 19456 37884 19508
rect 31760 19388 31812 19440
rect 33324 19431 33376 19440
rect 27068 19363 27120 19372
rect 27068 19329 27077 19363
rect 27077 19329 27111 19363
rect 27111 19329 27120 19363
rect 27068 19320 27120 19329
rect 27252 19363 27304 19372
rect 27252 19329 27261 19363
rect 27261 19329 27295 19363
rect 27295 19329 27304 19363
rect 27252 19320 27304 19329
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 32496 19363 32548 19372
rect 32496 19329 32505 19363
rect 32505 19329 32539 19363
rect 32539 19329 32548 19363
rect 32496 19320 32548 19329
rect 33324 19397 33358 19431
rect 33358 19397 33376 19431
rect 33324 19388 33376 19397
rect 33784 19388 33836 19440
rect 37188 19388 37240 19440
rect 40224 19388 40276 19440
rect 38752 19320 38804 19372
rect 39120 19363 39172 19372
rect 39120 19329 39129 19363
rect 39129 19329 39163 19363
rect 39163 19329 39172 19363
rect 39120 19320 39172 19329
rect 40316 19320 40368 19372
rect 40408 19320 40460 19372
rect 40776 19388 40828 19440
rect 41696 19431 41748 19440
rect 41696 19397 41705 19431
rect 41705 19397 41739 19431
rect 41739 19397 41748 19431
rect 46020 19456 46072 19508
rect 41696 19388 41748 19397
rect 40868 19363 40920 19372
rect 40868 19329 40877 19363
rect 40877 19329 40911 19363
rect 40911 19329 40920 19363
rect 40868 19320 40920 19329
rect 42616 19363 42668 19372
rect 42616 19329 42625 19363
rect 42625 19329 42659 19363
rect 42659 19329 42668 19363
rect 42616 19320 42668 19329
rect 43260 19363 43312 19372
rect 43260 19329 43269 19363
rect 43269 19329 43303 19363
rect 43303 19329 43312 19363
rect 43260 19320 43312 19329
rect 44640 19320 44692 19372
rect 45008 19363 45060 19372
rect 45008 19329 45022 19363
rect 45022 19329 45056 19363
rect 45056 19329 45060 19363
rect 45008 19320 45060 19329
rect 45192 19363 45244 19372
rect 45192 19329 45201 19363
rect 45201 19329 45235 19363
rect 45235 19329 45244 19363
rect 45192 19320 45244 19329
rect 46756 19320 46808 19372
rect 47768 19295 47820 19304
rect 41880 19227 41932 19236
rect 41880 19193 41889 19227
rect 41889 19193 41923 19227
rect 41923 19193 41932 19227
rect 41880 19184 41932 19193
rect 42064 19116 42116 19168
rect 47768 19261 47777 19295
rect 47777 19261 47811 19295
rect 47811 19261 47820 19295
rect 47768 19252 47820 19261
rect 45928 19116 45980 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 38844 18912 38896 18964
rect 40776 18912 40828 18964
rect 42064 18955 42116 18964
rect 42064 18921 42073 18955
rect 42073 18921 42107 18955
rect 42107 18921 42116 18955
rect 42064 18912 42116 18921
rect 42340 18912 42392 18964
rect 43536 18955 43588 18964
rect 38752 18887 38804 18896
rect 38752 18853 38761 18887
rect 38761 18853 38795 18887
rect 38795 18853 38804 18887
rect 38752 18844 38804 18853
rect 40040 18844 40092 18896
rect 43536 18921 43545 18955
rect 43545 18921 43579 18955
rect 43579 18921 43588 18955
rect 43536 18912 43588 18921
rect 44640 18912 44692 18964
rect 2136 18708 2188 18760
rect 2872 18708 2924 18760
rect 41604 18776 41656 18828
rect 40408 18751 40460 18760
rect 40408 18717 40417 18751
rect 40417 18717 40451 18751
rect 40451 18717 40460 18751
rect 40408 18708 40460 18717
rect 39212 18640 39264 18692
rect 2320 18572 2372 18624
rect 42064 18708 42116 18760
rect 42616 18708 42668 18760
rect 44364 18844 44416 18896
rect 45468 18844 45520 18896
rect 43628 18819 43680 18828
rect 43628 18785 43637 18819
rect 43637 18785 43671 18819
rect 43671 18785 43680 18819
rect 43628 18776 43680 18785
rect 46020 18776 46072 18828
rect 48136 18819 48188 18828
rect 48136 18785 48145 18819
rect 48145 18785 48179 18819
rect 48179 18785 48188 18819
rect 48136 18776 48188 18785
rect 44272 18751 44324 18760
rect 44272 18717 44281 18751
rect 44281 18717 44315 18751
rect 44315 18717 44324 18751
rect 44272 18708 44324 18717
rect 46296 18751 46348 18760
rect 46296 18717 46305 18751
rect 46305 18717 46339 18751
rect 46339 18717 46348 18751
rect 46296 18708 46348 18717
rect 43076 18640 43128 18692
rect 44088 18683 44140 18692
rect 44088 18649 44097 18683
rect 44097 18649 44131 18683
rect 44131 18649 44140 18683
rect 44088 18640 44140 18649
rect 46940 18640 46992 18692
rect 43168 18615 43220 18624
rect 43168 18581 43177 18615
rect 43177 18581 43211 18615
rect 43211 18581 43220 18615
rect 43168 18572 43220 18581
rect 44732 18572 44784 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 44456 18368 44508 18420
rect 45008 18411 45060 18420
rect 45008 18377 45017 18411
rect 45017 18377 45051 18411
rect 45051 18377 45060 18411
rect 45008 18368 45060 18377
rect 46940 18411 46992 18420
rect 46940 18377 46949 18411
rect 46949 18377 46983 18411
rect 46983 18377 46992 18411
rect 46940 18368 46992 18377
rect 2320 18343 2372 18352
rect 2320 18309 2329 18343
rect 2329 18309 2363 18343
rect 2363 18309 2372 18343
rect 2320 18300 2372 18309
rect 42616 18300 42668 18352
rect 42984 18300 43036 18352
rect 44180 18300 44232 18352
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 13636 18207 13688 18216
rect 13636 18173 13645 18207
rect 13645 18173 13679 18207
rect 13679 18173 13688 18207
rect 13636 18164 13688 18173
rect 15108 18207 15160 18216
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 42432 18164 42484 18216
rect 43536 18275 43588 18284
rect 43536 18241 43545 18275
rect 43545 18241 43579 18275
rect 43579 18241 43588 18275
rect 43536 18232 43588 18241
rect 44732 18275 44784 18284
rect 44732 18241 44741 18275
rect 44741 18241 44775 18275
rect 44775 18241 44784 18275
rect 44732 18232 44784 18241
rect 46296 18300 46348 18352
rect 46020 18232 46072 18284
rect 45468 18164 45520 18216
rect 47860 18164 47912 18216
rect 44088 18096 44140 18148
rect 42892 18028 42944 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 13636 17824 13688 17876
rect 15108 17824 15160 17876
rect 45560 17824 45612 17876
rect 39212 17799 39264 17808
rect 39212 17765 39221 17799
rect 39221 17765 39255 17799
rect 39255 17765 39264 17799
rect 39212 17756 39264 17765
rect 2136 17620 2188 17672
rect 12532 17620 12584 17672
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 37832 17663 37884 17672
rect 37832 17629 37841 17663
rect 37841 17629 37875 17663
rect 37875 17629 37884 17663
rect 37832 17620 37884 17629
rect 39856 17620 39908 17672
rect 42432 17756 42484 17808
rect 40500 17688 40552 17740
rect 42708 17756 42760 17808
rect 43076 17799 43128 17808
rect 43076 17765 43085 17799
rect 43085 17765 43119 17799
rect 43119 17765 43128 17799
rect 43076 17756 43128 17765
rect 42892 17688 42944 17740
rect 43168 17688 43220 17740
rect 42984 17620 43036 17672
rect 40960 17552 41012 17604
rect 44272 17620 44324 17672
rect 41144 17484 41196 17536
rect 41236 17484 41288 17536
rect 44088 17552 44140 17604
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 40408 17280 40460 17332
rect 44180 17323 44232 17332
rect 44180 17289 44189 17323
rect 44189 17289 44223 17323
rect 44223 17289 44232 17323
rect 44180 17280 44232 17289
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 40960 17187 41012 17196
rect 2320 17119 2372 17128
rect 2320 17085 2329 17119
rect 2329 17085 2363 17119
rect 2363 17085 2372 17119
rect 2320 17076 2372 17085
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 2780 17076 2832 17085
rect 40960 17153 40969 17187
rect 40969 17153 41003 17187
rect 41003 17153 41012 17187
rect 40960 17144 41012 17153
rect 41144 17187 41196 17196
rect 41144 17153 41153 17187
rect 41153 17153 41187 17187
rect 41187 17153 41196 17187
rect 41144 17144 41196 17153
rect 43628 17144 43680 17196
rect 44088 17187 44140 17196
rect 44088 17153 44097 17187
rect 44097 17153 44131 17187
rect 44131 17153 44140 17187
rect 44088 17144 44140 17153
rect 44272 17187 44324 17196
rect 44272 17153 44281 17187
rect 44281 17153 44315 17187
rect 44315 17153 44324 17187
rect 44272 17144 44324 17153
rect 47400 17144 47452 17196
rect 40224 17076 40276 17128
rect 42708 17119 42760 17128
rect 42708 17085 42717 17119
rect 42717 17085 42751 17119
rect 42751 17085 42760 17119
rect 42708 17076 42760 17085
rect 42984 17119 43036 17128
rect 42984 17085 42993 17119
rect 42993 17085 43027 17119
rect 43027 17085 43036 17119
rect 42984 17076 43036 17085
rect 40316 17008 40368 17060
rect 41236 17008 41288 17060
rect 46940 16983 46992 16992
rect 46940 16949 46949 16983
rect 46949 16949 46983 16983
rect 46983 16949 46992 16983
rect 46940 16940 46992 16949
rect 47768 16983 47820 16992
rect 47768 16949 47777 16983
rect 47777 16949 47811 16983
rect 47811 16949 47820 16983
rect 47768 16940 47820 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2320 16736 2372 16788
rect 39856 16779 39908 16788
rect 39856 16745 39865 16779
rect 39865 16745 39899 16779
rect 39899 16745 39908 16779
rect 39856 16736 39908 16745
rect 2412 16585 2464 16594
rect 2412 16551 2421 16585
rect 2421 16551 2455 16585
rect 2455 16551 2464 16585
rect 2412 16542 2464 16551
rect 40960 16600 41012 16652
rect 47768 16600 47820 16652
rect 48136 16643 48188 16652
rect 48136 16609 48145 16643
rect 48145 16609 48179 16643
rect 48179 16609 48188 16643
rect 48136 16600 48188 16609
rect 40408 16532 40460 16584
rect 46940 16464 46992 16516
rect 40224 16439 40276 16448
rect 40224 16405 40233 16439
rect 40233 16405 40267 16439
rect 40267 16405 40276 16439
rect 40224 16396 40276 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2136 15444 2188 15496
rect 47676 15487 47728 15496
rect 47676 15453 47685 15487
rect 47685 15453 47719 15487
rect 47719 15453 47728 15487
rect 47676 15444 47728 15453
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 47584 15011 47636 15020
rect 47584 14977 47593 15011
rect 47593 14977 47627 15011
rect 47627 14977 47636 15011
rect 47584 14968 47636 14977
rect 2596 14900 2648 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 46480 14764 46532 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2596 14603 2648 14612
rect 2596 14569 2605 14603
rect 2605 14569 2639 14603
rect 2639 14569 2648 14603
rect 2596 14560 2648 14569
rect 8576 14424 8628 14476
rect 9220 14424 9272 14476
rect 47676 14492 47728 14544
rect 46480 14467 46532 14476
rect 46480 14433 46489 14467
rect 46489 14433 46523 14467
rect 46523 14433 46532 14467
rect 46480 14424 46532 14433
rect 48136 14467 48188 14476
rect 48136 14433 48145 14467
rect 48145 14433 48179 14467
rect 48179 14433 48188 14467
rect 48136 14424 48188 14433
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 2136 14288 2188 14340
rect 2320 14220 2372 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2320 13991 2372 14000
rect 2320 13957 2329 13991
rect 2329 13957 2363 13991
rect 2363 13957 2372 13991
rect 2320 13948 2372 13957
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 46664 13744 46716 13796
rect 47124 13744 47176 13796
rect 47768 13719 47820 13728
rect 47768 13685 47777 13719
rect 47777 13685 47811 13719
rect 47811 13685 47820 13719
rect 47768 13676 47820 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 47768 13336 47820 13388
rect 48136 13379 48188 13388
rect 48136 13345 48145 13379
rect 48145 13345 48179 13379
rect 48179 13345 48188 13379
rect 48136 13336 48188 13345
rect 47676 13200 47728 13252
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 47676 12971 47728 12980
rect 47676 12937 47685 12971
rect 47685 12937 47719 12971
rect 47719 12937 47728 12971
rect 47676 12928 47728 12937
rect 46664 12792 46716 12844
rect 47584 12835 47636 12844
rect 47584 12801 47593 12835
rect 47593 12801 47627 12835
rect 47627 12801 47636 12835
rect 47584 12792 47636 12801
rect 46480 12588 46532 12640
rect 47032 12631 47084 12640
rect 47032 12597 47041 12631
rect 47041 12597 47075 12631
rect 47075 12597 47084 12631
rect 47032 12588 47084 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 47032 12316 47084 12368
rect 46480 12291 46532 12300
rect 46480 12257 46489 12291
rect 46489 12257 46523 12291
rect 46523 12257 46532 12291
rect 46480 12248 46532 12257
rect 48136 12291 48188 12300
rect 48136 12257 48145 12291
rect 48145 12257 48179 12291
rect 48179 12257 48188 12291
rect 48136 12248 48188 12257
rect 2044 12180 2096 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 18420 11704 18472 11756
rect 41420 11704 41472 11756
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 46480 11500 46532 11552
rect 47768 11543 47820 11552
rect 47768 11509 47777 11543
rect 47777 11509 47811 11543
rect 47811 11509 47820 11543
rect 47768 11500 47820 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2228 11296 2280 11348
rect 47768 11228 47820 11280
rect 46480 11203 46532 11212
rect 46480 11169 46489 11203
rect 46489 11169 46523 11203
rect 46523 11169 46532 11203
rect 46480 11160 46532 11169
rect 46848 11203 46900 11212
rect 46848 11169 46857 11203
rect 46857 11169 46891 11203
rect 46891 11169 46900 11203
rect 46848 11160 46900 11169
rect 2872 11092 2924 11144
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3148 10684 3200 10736
rect 2320 10591 2372 10600
rect 2320 10557 2329 10591
rect 2329 10557 2363 10591
rect 2363 10557 2372 10591
rect 2320 10548 2372 10557
rect 3700 10591 3752 10600
rect 3700 10557 3709 10591
rect 3709 10557 3743 10591
rect 3743 10557 3752 10591
rect 3700 10548 3752 10557
rect 5448 10412 5500 10464
rect 22100 10412 22152 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2320 10208 2372 10260
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 2780 10004 2832 10056
rect 5448 10004 5500 10056
rect 19984 10004 20036 10056
rect 20076 9979 20128 9988
rect 20076 9945 20085 9979
rect 20085 9945 20119 9979
rect 20119 9945 20128 9979
rect 20076 9936 20128 9945
rect 2964 9868 3016 9920
rect 27160 9868 27212 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2964 9639 3016 9648
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2780 9528 2832 9537
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 7196 9392 7248 9444
rect 2320 9324 2372 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2136 8916 2188 8968
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 45836 8576 45888 8628
rect 2320 8551 2372 8560
rect 2320 8517 2329 8551
rect 2329 8517 2363 8551
rect 2363 8517 2372 8551
rect 2320 8508 2372 8517
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 47952 8483 48004 8492
rect 47952 8449 47961 8483
rect 47961 8449 47995 8483
rect 47995 8449 48004 8483
rect 47952 8440 48004 8449
rect 2872 8415 2924 8424
rect 2872 8381 2881 8415
rect 2881 8381 2915 8415
rect 2915 8381 2924 8415
rect 2872 8372 2924 8381
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2228 7896 2280 7948
rect 2136 7828 2188 7880
rect 2964 7828 3016 7880
rect 2320 7692 2372 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2320 7463 2372 7472
rect 2320 7429 2329 7463
rect 2329 7429 2363 7463
rect 2363 7429 2372 7463
rect 2320 7420 2372 7429
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 47584 7395 47636 7404
rect 47584 7361 47593 7395
rect 47593 7361 47627 7395
rect 47627 7361 47636 7395
rect 47584 7352 47636 7361
rect 2780 7327 2832 7336
rect 2780 7293 2789 7327
rect 2789 7293 2823 7327
rect 2823 7293 2832 7327
rect 2780 7284 2832 7293
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 47676 7191 47728 7200
rect 47676 7157 47685 7191
rect 47685 7157 47719 7191
rect 47719 7157 47728 7191
rect 47676 7148 47728 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 47676 6808 47728 6860
rect 48136 6851 48188 6860
rect 48136 6817 48145 6851
rect 48145 6817 48179 6851
rect 48179 6817 48188 6851
rect 48136 6808 48188 6817
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 47768 6672 47820 6724
rect 2320 6604 2372 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2320 6375 2372 6384
rect 2320 6341 2329 6375
rect 2329 6341 2363 6375
rect 2363 6341 2372 6375
rect 2320 6332 2372 6341
rect 1676 6264 1728 6316
rect 45560 6264 45612 6316
rect 47492 6332 47544 6384
rect 46664 6264 46716 6316
rect 47768 6307 47820 6316
rect 47768 6273 47777 6307
rect 47777 6273 47811 6307
rect 47811 6273 47820 6307
rect 47768 6264 47820 6273
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 46296 6103 46348 6112
rect 46296 6069 46305 6103
rect 46305 6069 46339 6103
rect 46339 6069 46348 6103
rect 46296 6060 46348 6069
rect 46940 6103 46992 6112
rect 46940 6069 46949 6103
rect 46949 6069 46983 6103
rect 46983 6069 46992 6103
rect 46940 6060 46992 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1676 5652 1728 5704
rect 2412 5652 2464 5704
rect 17224 5652 17276 5704
rect 17868 5652 17920 5704
rect 45652 5695 45704 5704
rect 45652 5661 45661 5695
rect 45661 5661 45695 5695
rect 45695 5661 45704 5695
rect 45652 5652 45704 5661
rect 45836 5652 45888 5704
rect 48228 5584 48280 5636
rect 3884 5559 3936 5568
rect 3884 5525 3893 5559
rect 3893 5525 3927 5559
rect 3927 5525 3936 5559
rect 3884 5516 3936 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2780 5312 2832 5364
rect 4068 5312 4120 5364
rect 3884 5244 3936 5296
rect 46296 5244 46348 5296
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 46848 5151 46900 5160
rect 46848 5117 46857 5151
rect 46857 5117 46891 5151
rect 46891 5117 46900 5151
rect 46848 5108 46900 5117
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 46296 4972 46348 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2872 4632 2924 4684
rect 2780 4564 2832 4616
rect 8024 4768 8076 4820
rect 14096 4768 14148 4820
rect 45836 4768 45888 4820
rect 46296 4675 46348 4684
rect 46296 4641 46305 4675
rect 46305 4641 46339 4675
rect 46339 4641 46348 4675
rect 46296 4632 46348 4641
rect 46940 4632 46992 4684
rect 48136 4675 48188 4684
rect 48136 4641 48145 4675
rect 48145 4641 48179 4675
rect 48179 4641 48188 4675
rect 48136 4632 48188 4641
rect 4712 4564 4764 4616
rect 3976 4496 4028 4548
rect 4528 4496 4580 4548
rect 6092 4564 6144 4616
rect 7748 4564 7800 4616
rect 9036 4564 9088 4616
rect 17316 4564 17368 4616
rect 20076 4564 20128 4616
rect 42340 4607 42392 4616
rect 42340 4573 42349 4607
rect 42349 4573 42383 4607
rect 42383 4573 42392 4607
rect 42340 4564 42392 4573
rect 46204 4564 46256 4616
rect 20444 4496 20496 4548
rect 2412 4471 2464 4480
rect 2412 4437 2421 4471
rect 2421 4437 2455 4471
rect 2455 4437 2464 4471
rect 2412 4428 2464 4437
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 4988 4471 5040 4480
rect 4988 4437 4997 4471
rect 4997 4437 5031 4471
rect 5031 4437 5040 4471
rect 4988 4428 5040 4437
rect 8576 4428 8628 4480
rect 19340 4471 19392 4480
rect 19340 4437 19349 4471
rect 19349 4437 19383 4471
rect 19383 4437 19392 4471
rect 19340 4428 19392 4437
rect 19984 4471 20036 4480
rect 19984 4437 19993 4471
rect 19993 4437 20027 4471
rect 20027 4437 20036 4471
rect 19984 4428 20036 4437
rect 45376 4471 45428 4480
rect 45376 4437 45385 4471
rect 45385 4437 45419 4471
rect 45419 4437 45428 4471
rect 45376 4428 45428 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 1492 4131 1544 4140
rect 1492 4097 1501 4131
rect 1501 4097 1535 4131
rect 1535 4097 1544 4131
rect 1492 4088 1544 4097
rect 1952 4088 2004 4140
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 7196 4088 7248 4140
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 38660 4131 38712 4140
rect 3056 4020 3108 4072
rect 3148 4063 3200 4072
rect 3148 4029 3157 4063
rect 3157 4029 3191 4063
rect 3191 4029 3200 4063
rect 3148 4020 3200 4029
rect 8576 4020 8628 4072
rect 12348 4063 12400 4072
rect 7104 3952 7156 4004
rect 12348 4029 12357 4063
rect 12357 4029 12391 4063
rect 12391 4029 12400 4063
rect 12348 4020 12400 4029
rect 12808 4020 12860 4072
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 19340 4020 19392 4072
rect 19432 4063 19484 4072
rect 19432 4029 19441 4063
rect 19441 4029 19475 4063
rect 19475 4029 19484 4063
rect 19432 4020 19484 4029
rect 9220 3952 9272 4004
rect 38660 4097 38669 4131
rect 38669 4097 38703 4131
rect 38703 4097 38712 4131
rect 41512 4224 41564 4276
rect 38660 4088 38712 4097
rect 38568 3952 38620 4004
rect 41972 4156 42024 4208
rect 40776 4131 40828 4140
rect 40776 4097 40785 4131
rect 40785 4097 40819 4131
rect 40819 4097 40828 4131
rect 40776 4088 40828 4097
rect 42524 4088 42576 4140
rect 45560 4224 45612 4276
rect 45376 4199 45428 4208
rect 45376 4165 45385 4199
rect 45385 4165 45419 4199
rect 45419 4165 45428 4199
rect 45376 4156 45428 4165
rect 47032 4063 47084 4072
rect 41420 3952 41472 4004
rect 41512 3952 41564 4004
rect 47032 4029 47041 4063
rect 47041 4029 47075 4063
rect 47075 4029 47084 4063
rect 47032 4020 47084 4029
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 6276 3884 6328 3936
rect 9128 3884 9180 3936
rect 10416 3884 10468 3936
rect 17132 3884 17184 3936
rect 22192 3927 22244 3936
rect 22192 3893 22201 3927
rect 22201 3893 22235 3927
rect 22235 3893 22244 3927
rect 22192 3884 22244 3893
rect 25504 3927 25556 3936
rect 25504 3893 25513 3927
rect 25513 3893 25547 3927
rect 25547 3893 25556 3927
rect 25504 3884 25556 3893
rect 38752 3927 38804 3936
rect 38752 3893 38761 3927
rect 38761 3893 38795 3927
rect 38795 3893 38804 3927
rect 38752 3884 38804 3893
rect 40040 3884 40092 3936
rect 40868 3927 40920 3936
rect 40868 3893 40877 3927
rect 40877 3893 40911 3927
rect 40911 3893 40920 3927
rect 40868 3884 40920 3893
rect 41788 3927 41840 3936
rect 41788 3893 41797 3927
rect 41797 3893 41831 3927
rect 41831 3893 41840 3927
rect 41788 3884 41840 3893
rect 42156 3884 42208 3936
rect 43628 3927 43680 3936
rect 43628 3893 43637 3927
rect 43637 3893 43671 3927
rect 43671 3893 43680 3927
rect 43628 3884 43680 3893
rect 44732 3884 44784 3936
rect 47584 3884 47636 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 14096 3680 14148 3732
rect 1492 3612 1544 3664
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 3976 3587 4028 3596
rect 3976 3553 3985 3587
rect 3985 3553 4019 3587
rect 4019 3553 4028 3587
rect 3976 3544 4028 3553
rect 4068 3544 4120 3596
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 6460 3544 6512 3596
rect 7196 3612 7248 3664
rect 9404 3544 9456 3596
rect 10416 3587 10468 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 9680 3476 9732 3528
rect 7840 3408 7892 3460
rect 8024 3340 8076 3392
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 17868 3612 17920 3664
rect 25596 3612 25648 3664
rect 10692 3408 10744 3460
rect 13452 3476 13504 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 20076 3544 20128 3596
rect 25504 3587 25556 3596
rect 25504 3553 25513 3587
rect 25513 3553 25547 3587
rect 25547 3553 25556 3587
rect 25504 3544 25556 3553
rect 25780 3680 25832 3732
rect 28172 3612 28224 3664
rect 41880 3680 41932 3732
rect 28356 3612 28408 3664
rect 40040 3587 40092 3596
rect 13636 3340 13688 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 22008 3476 22060 3528
rect 25320 3519 25372 3528
rect 25320 3485 25329 3519
rect 25329 3485 25363 3519
rect 25363 3485 25372 3519
rect 25320 3476 25372 3485
rect 21364 3451 21416 3460
rect 21364 3417 21373 3451
rect 21373 3417 21407 3451
rect 21407 3417 21416 3451
rect 21364 3408 21416 3417
rect 25780 3408 25832 3460
rect 27804 3519 27856 3528
rect 27804 3485 27813 3519
rect 27813 3485 27847 3519
rect 27847 3485 27856 3519
rect 27804 3476 27856 3485
rect 32128 3476 32180 3528
rect 40040 3553 40049 3587
rect 40049 3553 40083 3587
rect 40083 3553 40092 3587
rect 40040 3544 40092 3553
rect 40592 3587 40644 3596
rect 40592 3553 40601 3587
rect 40601 3553 40635 3587
rect 40635 3553 40644 3587
rect 40592 3544 40644 3553
rect 41788 3612 41840 3664
rect 41972 3544 42024 3596
rect 42156 3587 42208 3596
rect 42156 3553 42165 3587
rect 42165 3553 42199 3587
rect 42199 3553 42208 3587
rect 42156 3544 42208 3553
rect 18604 3340 18656 3392
rect 28356 3383 28408 3392
rect 28356 3349 28365 3383
rect 28365 3349 28399 3383
rect 28399 3349 28408 3383
rect 28356 3340 28408 3349
rect 32312 3383 32364 3392
rect 32312 3349 32321 3383
rect 32321 3349 32355 3383
rect 32355 3349 32364 3383
rect 32312 3340 32364 3349
rect 38476 3408 38528 3460
rect 43352 3408 43404 3460
rect 45652 3680 45704 3732
rect 46388 3612 46440 3664
rect 47492 3544 47544 3596
rect 47768 3587 47820 3596
rect 47768 3553 47777 3587
rect 47777 3553 47811 3587
rect 47811 3553 47820 3587
rect 47768 3544 47820 3553
rect 45836 3519 45888 3528
rect 45836 3485 45845 3519
rect 45845 3485 45879 3519
rect 45879 3485 45888 3519
rect 45836 3476 45888 3485
rect 47676 3408 47728 3460
rect 45192 3340 45244 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 10692 3179 10744 3188
rect 2412 3068 2464 3120
rect 4620 3068 4672 3120
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 8024 3111 8076 3120
rect 8024 3077 8033 3111
rect 8033 3077 8067 3111
rect 8067 3077 8076 3111
rect 8024 3068 8076 3077
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 9680 3068 9732 3120
rect 18880 3136 18932 3188
rect 13636 3111 13688 3120
rect 13636 3077 13645 3111
rect 13645 3077 13679 3111
rect 13679 3077 13688 3111
rect 13636 3068 13688 3077
rect 17316 3111 17368 3120
rect 17316 3077 17325 3111
rect 17325 3077 17359 3111
rect 17359 3077 17368 3111
rect 17316 3068 17368 3077
rect 19984 3068 20036 3120
rect 21364 3136 21416 3188
rect 38476 3136 38528 3188
rect 47676 3179 47728 3188
rect 38752 3111 38804 3120
rect 38752 3077 38761 3111
rect 38761 3077 38795 3111
rect 38795 3077 38804 3111
rect 38752 3068 38804 3077
rect 40868 3068 40920 3120
rect 47676 3145 47685 3179
rect 47685 3145 47719 3179
rect 47719 3145 47728 3179
rect 47676 3136 47728 3145
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 4712 2932 4764 2984
rect 12348 3000 12400 3052
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 25320 3000 25372 3052
rect 32128 3043 32180 3052
rect 32128 3009 32137 3043
rect 32137 3009 32171 3043
rect 32171 3009 32180 3043
rect 32128 3000 32180 3009
rect 38568 3043 38620 3052
rect 38568 3009 38577 3043
rect 38577 3009 38611 3043
rect 38611 3009 38620 3043
rect 38568 3000 38620 3009
rect 664 2864 716 2916
rect 5172 2864 5224 2916
rect 13084 2932 13136 2984
rect 17408 2932 17460 2984
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 22192 2975 22244 2984
rect 22192 2941 22201 2975
rect 22201 2941 22235 2975
rect 22235 2941 22244 2975
rect 22192 2932 22244 2941
rect 22560 2975 22612 2984
rect 22560 2941 22569 2975
rect 22569 2941 22603 2975
rect 22603 2941 22612 2975
rect 22560 2932 22612 2941
rect 27160 2975 27212 2984
rect 27160 2941 27169 2975
rect 27169 2941 27203 2975
rect 27203 2941 27212 2975
rect 27160 2932 27212 2941
rect 27252 2932 27304 2984
rect 32312 2975 32364 2984
rect 32312 2941 32321 2975
rect 32321 2941 32355 2975
rect 32355 2941 32364 2975
rect 32312 2932 32364 2941
rect 32404 2932 32456 2984
rect 39304 2975 39356 2984
rect 39304 2941 39313 2975
rect 39313 2941 39347 2975
rect 39347 2941 39356 2975
rect 39304 2932 39356 2941
rect 13544 2864 13596 2916
rect 6552 2796 6604 2848
rect 8944 2796 8996 2848
rect 9496 2796 9548 2848
rect 38660 2864 38712 2916
rect 18788 2796 18840 2848
rect 40776 3000 40828 3052
rect 44732 3043 44784 3052
rect 44732 3009 44741 3043
rect 44741 3009 44775 3043
rect 44775 3009 44784 3043
rect 44732 3000 44784 3009
rect 41236 2864 41288 2916
rect 43628 2932 43680 2984
rect 46572 2975 46624 2984
rect 46572 2941 46581 2975
rect 46581 2941 46615 2975
rect 46615 2941 46624 2975
rect 46572 2932 46624 2941
rect 43352 2864 43404 2916
rect 45744 2864 45796 2916
rect 42616 2796 42668 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1400 2592 1452 2644
rect 19432 2592 19484 2644
rect 47492 2592 47544 2644
rect 3792 2524 3844 2576
rect 4528 2524 4580 2576
rect 3332 2456 3384 2508
rect 5816 2456 5868 2508
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 7748 2524 7800 2576
rect 8944 2499 8996 2508
rect 8944 2465 8953 2499
rect 8953 2465 8987 2499
rect 8987 2465 8996 2499
rect 8944 2456 8996 2465
rect 9128 2499 9180 2508
rect 9128 2465 9137 2499
rect 9137 2465 9171 2499
rect 9171 2465 9180 2499
rect 9128 2456 9180 2465
rect 24216 2456 24268 2508
rect 27804 2524 27856 2576
rect 28356 2456 28408 2508
rect 23848 2388 23900 2440
rect 4988 2320 5040 2372
rect 27712 2320 27764 2372
rect 42340 2456 42392 2508
rect 42616 2499 42668 2508
rect 42616 2465 42625 2499
rect 42625 2465 42659 2499
rect 42659 2465 42668 2499
rect 42616 2456 42668 2465
rect 45836 2524 45888 2576
rect 45192 2499 45244 2508
rect 45192 2465 45201 2499
rect 45201 2465 45235 2499
rect 45235 2465 45244 2499
rect 45192 2456 45244 2465
rect 45284 2456 45336 2508
rect 48964 2320 49016 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect -10 49200 102 50000
rect 1278 49200 1390 50000
rect 1922 49314 2034 50000
rect 1922 49286 2176 49314
rect 1922 49200 2034 49286
rect 32 47122 60 49200
rect 20 47116 72 47122
rect 20 47058 72 47064
rect 2148 46510 2176 49286
rect 2566 49200 2678 50000
rect 3854 49200 3966 50000
rect 4498 49200 4610 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7718 49200 7830 50000
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 10294 49200 10406 50000
rect 10938 49200 11050 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18666 49200 18778 50000
rect 19310 49200 19422 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 21886 49200 21998 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 25106 49200 25218 50000
rect 25750 49200 25862 50000
rect 27038 49200 27150 50000
rect 27682 49314 27794 50000
rect 27682 49286 28028 49314
rect 27682 49200 27794 49286
rect 2608 46714 2636 49200
rect 3606 48376 3662 48385
rect 3606 48311 3662 48320
rect 2778 47696 2834 47705
rect 2778 47631 2834 47640
rect 2688 47048 2740 47054
rect 2688 46990 2740 46996
rect 2596 46708 2648 46714
rect 2596 46650 2648 46656
rect 2136 46504 2188 46510
rect 2136 46446 2188 46452
rect 1768 46436 1820 46442
rect 1768 46378 1820 46384
rect 1674 46336 1730 46345
rect 1674 46271 1730 46280
rect 1400 45960 1452 45966
rect 1400 45902 1452 45908
rect 1412 45082 1440 45902
rect 1688 45558 1716 46271
rect 1676 45552 1728 45558
rect 1676 45494 1728 45500
rect 1400 45076 1452 45082
rect 1400 45018 1452 45024
rect 1780 45014 1808 46378
rect 1768 45008 1820 45014
rect 1768 44950 1820 44956
rect 2136 43784 2188 43790
rect 2136 43726 2188 43732
rect 2148 43314 2176 43726
rect 2136 43308 2188 43314
rect 2136 43250 2188 43256
rect 2700 40594 2728 46990
rect 2792 46034 2820 47631
rect 2964 47184 3016 47190
rect 2964 47126 3016 47132
rect 2872 46980 2924 46986
rect 2872 46922 2924 46928
rect 2780 46028 2832 46034
rect 2780 45970 2832 45976
rect 2884 45558 2912 46922
rect 2872 45552 2924 45558
rect 2872 45494 2924 45500
rect 2976 45422 3004 47126
rect 3056 46708 3108 46714
rect 3056 46650 3108 46656
rect 3068 45422 3096 46650
rect 3148 45892 3200 45898
rect 3148 45834 3200 45840
rect 2964 45416 3016 45422
rect 2964 45358 3016 45364
rect 3056 45416 3108 45422
rect 3056 45358 3108 45364
rect 3160 45082 3188 45834
rect 3148 45076 3200 45082
rect 3148 45018 3200 45024
rect 3056 44872 3108 44878
rect 3056 44814 3108 44820
rect 3068 44538 3096 44814
rect 3056 44532 3108 44538
rect 3056 44474 3108 44480
rect 2688 40588 2740 40594
rect 2688 40530 2740 40536
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 2056 34610 2084 35022
rect 2044 34604 2096 34610
rect 2044 34546 2096 34552
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 2240 34202 2268 34478
rect 2228 34196 2280 34202
rect 2228 34138 2280 34144
rect 2412 33992 2464 33998
rect 2412 33934 2464 33940
rect 2136 32904 2188 32910
rect 2136 32846 2188 32852
rect 2148 32434 2176 32846
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 2424 26234 2452 33934
rect 2778 32736 2834 32745
rect 2778 32671 2834 32680
rect 2792 32366 2820 32671
rect 2504 32360 2556 32366
rect 2504 32302 2556 32308
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2516 32026 2544 32302
rect 2504 32020 2556 32026
rect 2504 31962 2556 31968
rect 2424 26206 2544 26234
rect 2136 25288 2188 25294
rect 2136 25230 2188 25236
rect 2148 24818 2176 25230
rect 2320 25152 2372 25158
rect 2320 25094 2372 25100
rect 2332 24886 2360 25094
rect 2320 24880 2372 24886
rect 2320 24822 2372 24828
rect 2136 24812 2188 24818
rect 2136 24754 2188 24760
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 2056 23730 2084 24142
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 2228 23656 2280 23662
rect 2228 23598 2280 23604
rect 2240 23322 2268 23598
rect 2228 23316 2280 23322
rect 2228 23258 2280 23264
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2044 22024 2096 22030
rect 2044 21966 2096 21972
rect 2056 21554 2084 21966
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2148 18290 2176 18702
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2148 17202 2176 17614
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2148 15026 2176 15438
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2148 13938 2176 14282
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 11762 2084 12174
rect 2240 11778 2268 23054
rect 2412 21480 2464 21486
rect 2412 21422 2464 21428
rect 2424 21146 2452 21422
rect 2412 21140 2464 21146
rect 2412 21082 2464 21088
rect 2516 19802 2544 26206
rect 3068 25770 3096 44474
rect 3330 41576 3386 41585
rect 3330 41511 3386 41520
rect 3344 35894 3372 41511
rect 3424 40996 3476 41002
rect 3424 40938 3476 40944
rect 3436 40905 3464 40938
rect 3422 40896 3478 40905
rect 3422 40831 3478 40840
rect 3344 35866 3464 35894
rect 3056 25764 3108 25770
rect 3056 25706 3108 25712
rect 2778 25256 2834 25265
rect 2778 25191 2834 25200
rect 2792 24750 2820 25191
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 3436 24682 3464 35866
rect 3620 34542 3648 48311
rect 4540 47954 4568 49200
rect 4540 47926 4660 47954
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4252 47048 4304 47054
rect 4252 46990 4304 46996
rect 4264 46646 4292 46990
rect 3884 46640 3936 46646
rect 3884 46582 3936 46588
rect 4252 46640 4304 46646
rect 4252 46582 4304 46588
rect 3698 45656 3754 45665
rect 3698 45591 3754 45600
rect 3608 34536 3660 34542
rect 3608 34478 3660 34484
rect 3424 24676 3476 24682
rect 3424 24618 3476 24624
rect 2778 23896 2834 23905
rect 2778 23831 2834 23840
rect 2792 23662 2820 23831
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2778 21856 2834 21865
rect 2778 21791 2834 21800
rect 2792 21486 2820 21791
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2884 20942 2912 21354
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 2778 20496 2834 20505
rect 2778 20431 2834 20440
rect 2792 20398 2820 20431
rect 2596 20392 2648 20398
rect 2596 20334 2648 20340
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2608 20058 2636 20334
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2424 19774 2544 19802
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2332 18358 2360 18566
rect 2320 18352 2372 18358
rect 2320 18294 2372 18300
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 2332 16794 2360 17070
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2424 16600 2452 19774
rect 2504 19712 2556 19718
rect 2504 19654 2556 19660
rect 2412 16594 2464 16600
rect 2412 16536 2464 16542
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2332 14006 2360 14214
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2148 11750 2268 11778
rect 2148 10146 2176 11750
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11354 2268 11630
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 10266 2360 10542
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2148 10118 2268 10146
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 9586 2176 9998
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8498 2176 8910
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2240 7954 2268 10118
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 8566 2360 9318
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 7410 2176 7822
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2332 7478 2360 7686
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6322 1716 7142
rect 2424 6798 2452 16536
rect 2516 14414 2544 19654
rect 2884 18766 2912 20878
rect 3160 20534 3188 20878
rect 3148 20528 3200 20534
rect 3148 20470 3200 20476
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2792 18222 2820 18391
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 2780 17128 2832 17134
rect 2778 17096 2780 17105
rect 2832 17096 2834 17105
rect 2778 17031 2834 17040
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 14958 2820 14991
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2608 14618 2636 14894
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2778 14376 2834 14385
rect 2778 14311 2834 14320
rect 2792 13870 2820 14311
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2780 11688 2832 11694
rect 2778 11656 2780 11665
rect 2832 11656 2834 11665
rect 2778 11591 2834 11600
rect 2884 11150 2912 18702
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10742 3188 11086
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3712 10606 3740 45591
rect 3896 45082 3924 46582
rect 4632 46510 4660 47926
rect 5540 47048 5592 47054
rect 5540 46990 5592 46996
rect 4620 46504 4672 46510
rect 4620 46446 4672 46452
rect 4068 46436 4120 46442
rect 4068 46378 4120 46384
rect 4080 46170 4108 46378
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4068 46164 4120 46170
rect 4068 46106 4120 46112
rect 5552 46034 5580 46990
rect 5828 46034 5856 49200
rect 8404 47054 8432 49200
rect 8392 47048 8444 47054
rect 8392 46990 8444 46996
rect 8944 46912 8996 46918
rect 8944 46854 8996 46860
rect 5540 46028 5592 46034
rect 5540 45970 5592 45976
rect 5816 46028 5868 46034
rect 5816 45970 5868 45976
rect 5540 45892 5592 45898
rect 5540 45834 5592 45840
rect 4068 45824 4120 45830
rect 4068 45766 4120 45772
rect 3884 45076 3936 45082
rect 3884 45018 3936 45024
rect 3974 43616 4030 43625
rect 3974 43551 4030 43560
rect 3988 43382 4016 43551
rect 3976 43376 4028 43382
rect 3976 43318 4028 43324
rect 3884 43240 3936 43246
rect 3884 43182 3936 43188
rect 3896 42770 3924 43182
rect 3884 42764 3936 42770
rect 3884 42706 3936 42712
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3238 10296 3294 10305
rect 3238 10231 3294 10240
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2792 9586 2820 9998
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9654 3004 9862
rect 2964 9648 3016 9654
rect 2870 9616 2926 9625
rect 2780 9580 2832 9586
rect 2964 9590 3016 9596
rect 2870 9551 2926 9560
rect 2780 9522 2832 9528
rect 2884 8430 2912 9551
rect 3252 9518 3280 10231
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2778 7576 2834 7585
rect 2778 7511 2834 7520
rect 2792 7342 2820 7511
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 6390 2360 6598
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 2792 6254 2820 6831
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1504 3670 1532 4082
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1492 3664 1544 3670
rect 1492 3606 1544 3612
rect 1596 3602 1624 3878
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 664 2916 716 2922
rect 664 2858 716 2864
rect 676 800 704 2858
rect 1412 2650 1440 3470
rect 1688 3058 1716 5646
rect 2424 5234 2452 5646
rect 2870 5536 2926 5545
rect 2870 5471 2926 5480
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1964 4146 1992 4966
rect 2792 4622 2820 5306
rect 2884 5166 2912 5471
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2976 4978 3004 7822
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5302 3924 5510
rect 4080 5370 4108 45766
rect 5552 45558 5580 45834
rect 5540 45552 5592 45558
rect 5540 45494 5592 45500
rect 5448 45484 5500 45490
rect 5448 45426 5500 45432
rect 8392 45484 8444 45490
rect 8392 45426 8444 45432
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5460 10470 5488 45426
rect 8404 45354 8432 45426
rect 8392 45348 8444 45354
rect 8392 45290 8444 45296
rect 8208 44940 8260 44946
rect 8208 44882 8260 44888
rect 6368 42696 6420 42702
rect 6368 42638 6420 42644
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 5460 10062 5488 10406
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 2884 4950 3004 4978
rect 2884 4690 2912 4950
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 3146 4856 3202 4865
rect 4214 4859 4522 4868
rect 3146 4791 3202 4800
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3505 1900 3538
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 2424 3126 2452 4422
rect 3068 4078 3096 4422
rect 3160 4078 3188 4791
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3988 3602 4016 4490
rect 4540 4146 4568 4490
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 2792 1465 2820 2926
rect 3804 2582 3832 3470
rect 4080 2825 4108 3538
rect 4632 3126 4660 3878
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4724 2990 4752 4558
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4066 2816 4122 2825
rect 4066 2751 4122 2760
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3792 2576 3844 2582
rect 3792 2518 3844 2524
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3344 1170 3372 2450
rect 3252 1142 3372 1170
rect 3252 800 3280 1142
rect 4540 800 4568 2518
rect 5000 2378 5028 4422
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 5184 800 5212 2858
rect 5828 2514 5856 3878
rect 6104 3602 6132 4558
rect 6380 4146 6408 42638
rect 7932 26784 7984 26790
rect 7932 26726 7984 26732
rect 7944 26382 7972 26726
rect 8220 26586 8248 44882
rect 8404 27470 8432 45290
rect 8956 42634 8984 46854
rect 9588 46436 9640 46442
rect 9588 46378 9640 46384
rect 9600 46034 9628 46378
rect 10876 46368 10928 46374
rect 10876 46310 10928 46316
rect 10888 46034 10916 46310
rect 10980 46102 11008 49200
rect 11520 47116 11572 47122
rect 11520 47058 11572 47064
rect 10968 46096 11020 46102
rect 10968 46038 11020 46044
rect 9588 46028 9640 46034
rect 9588 45970 9640 45976
rect 10876 46028 10928 46034
rect 10876 45970 10928 45976
rect 9220 45960 9272 45966
rect 9220 45902 9272 45908
rect 9232 45490 9260 45902
rect 9600 45558 9628 45970
rect 10784 45824 10836 45830
rect 10784 45766 10836 45772
rect 9588 45552 9640 45558
rect 9588 45494 9640 45500
rect 9220 45484 9272 45490
rect 9220 45426 9272 45432
rect 9232 44878 9260 45426
rect 10796 45422 10824 45766
rect 11532 45490 11560 47058
rect 12716 47048 12768 47054
rect 12716 46990 12768 46996
rect 12728 46646 12756 46990
rect 12716 46640 12768 46646
rect 12716 46582 12768 46588
rect 12912 46510 12940 49200
rect 14200 47410 14228 49200
rect 14200 47382 14320 47410
rect 13176 47048 13228 47054
rect 13176 46990 13228 46996
rect 14188 47048 14240 47054
rect 14188 46990 14240 46996
rect 12624 46504 12676 46510
rect 12624 46446 12676 46452
rect 12900 46504 12952 46510
rect 12900 46446 12952 46452
rect 12532 45960 12584 45966
rect 12532 45902 12584 45908
rect 11612 45892 11664 45898
rect 11612 45834 11664 45840
rect 11624 45626 11652 45834
rect 11612 45620 11664 45626
rect 11612 45562 11664 45568
rect 12544 45490 12572 45902
rect 12636 45558 12664 46446
rect 12624 45552 12676 45558
rect 12624 45494 12676 45500
rect 13188 45490 13216 46990
rect 14200 46578 14228 46990
rect 14188 46572 14240 46578
rect 14188 46514 14240 46520
rect 13360 45824 13412 45830
rect 13360 45766 13412 45772
rect 13372 45558 13400 45766
rect 13360 45552 13412 45558
rect 13360 45494 13412 45500
rect 11520 45484 11572 45490
rect 11520 45426 11572 45432
rect 12532 45484 12584 45490
rect 12532 45426 12584 45432
rect 13176 45484 13228 45490
rect 13176 45426 13228 45432
rect 9404 45416 9456 45422
rect 9404 45358 9456 45364
rect 10784 45416 10836 45422
rect 10784 45358 10836 45364
rect 9416 45014 9444 45358
rect 9404 45008 9456 45014
rect 9404 44950 9456 44956
rect 9220 44872 9272 44878
rect 9220 44814 9272 44820
rect 9232 44402 9260 44814
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 9036 44328 9088 44334
rect 9036 44270 9088 44276
rect 8944 42628 8996 42634
rect 8944 42570 8996 42576
rect 8852 41064 8904 41070
rect 8852 41006 8904 41012
rect 8864 40730 8892 41006
rect 8852 40724 8904 40730
rect 8852 40666 8904 40672
rect 8576 31816 8628 31822
rect 8576 31758 8628 31764
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8404 27062 8432 27406
rect 8392 27056 8444 27062
rect 8392 26998 8444 27004
rect 8208 26580 8260 26586
rect 8208 26522 8260 26528
rect 8220 26450 8248 26522
rect 8208 26444 8260 26450
rect 8208 26386 8260 26392
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 7944 26234 7972 26318
rect 7852 26206 7972 26234
rect 7852 25906 7880 26206
rect 8588 25974 8616 31758
rect 8576 25968 8628 25974
rect 8576 25910 8628 25916
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7852 25294 7880 25842
rect 8588 25838 8616 25910
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 7852 24818 7880 25230
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 8024 24744 8076 24750
rect 8024 24686 8076 24692
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 4146 7236 9386
rect 8036 4826 8064 24686
rect 8588 14482 8616 25774
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 9048 4622 9076 44270
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 7760 4146 7788 4558
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6288 3602 6316 3878
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6472 800 6500 3538
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2514 6592 2790
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 7116 800 7144 3946
rect 7208 3670 7236 4082
rect 8588 4078 8616 4422
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 9232 4010 9260 14418
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7852 3058 7880 3402
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8036 3126 8064 3334
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7760 800 7788 2518
rect 8956 2514 8984 2790
rect 9140 2514 9168 3878
rect 9416 3602 9444 44950
rect 9588 44804 9640 44810
rect 9588 44746 9640 44752
rect 9600 42702 9628 44746
rect 9588 42696 9640 42702
rect 9588 42638 9640 42644
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9508 2854 9536 25774
rect 12544 25294 12572 45426
rect 14292 45422 14320 47382
rect 14844 46510 14872 49200
rect 14464 46504 14516 46510
rect 14464 46446 14516 46452
rect 14832 46504 14884 46510
rect 14832 46446 14884 46452
rect 14476 46170 14504 46446
rect 14464 46164 14516 46170
rect 14464 46106 14516 46112
rect 15488 46102 15516 49200
rect 15660 47048 15712 47054
rect 15660 46990 15712 46996
rect 15476 46096 15528 46102
rect 15476 46038 15528 46044
rect 15672 46034 15700 46990
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 23216 46510 23244 49200
rect 24860 47048 24912 47054
rect 24860 46990 24912 46996
rect 22284 46504 22336 46510
rect 22284 46446 22336 46452
rect 22928 46504 22980 46510
rect 22928 46446 22980 46452
rect 23204 46504 23256 46510
rect 23204 46446 23256 46452
rect 17224 46436 17276 46442
rect 17224 46378 17276 46384
rect 17236 46034 17264 46378
rect 22296 46170 22324 46446
rect 22284 46164 22336 46170
rect 22284 46106 22336 46112
rect 15660 46028 15712 46034
rect 15660 45970 15712 45976
rect 17224 46028 17276 46034
rect 17224 45970 17276 45976
rect 15568 45892 15620 45898
rect 15568 45834 15620 45840
rect 14372 45824 14424 45830
rect 14372 45766 14424 45772
rect 14280 45416 14332 45422
rect 14280 45358 14332 45364
rect 14384 44946 14412 45766
rect 15580 45626 15608 45834
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 22940 45626 22968 46446
rect 24872 46050 24900 46990
rect 24688 46022 24900 46050
rect 24688 45966 24716 46022
rect 24676 45960 24728 45966
rect 24676 45902 24728 45908
rect 25148 45898 25176 49200
rect 25504 47048 25556 47054
rect 25504 46990 25556 46996
rect 25516 46646 25544 46990
rect 25504 46640 25556 46646
rect 25504 46582 25556 46588
rect 25792 46510 25820 49200
rect 26424 47048 26476 47054
rect 26424 46990 26476 46996
rect 26436 46578 26464 46990
rect 26424 46572 26476 46578
rect 26424 46514 26476 46520
rect 25320 46504 25372 46510
rect 25320 46446 25372 46452
rect 25780 46504 25832 46510
rect 25780 46446 25832 46452
rect 26240 46504 26292 46510
rect 26240 46446 26292 46452
rect 24860 45892 24912 45898
rect 24860 45834 24912 45840
rect 25136 45892 25188 45898
rect 25136 45834 25188 45840
rect 15568 45620 15620 45626
rect 15568 45562 15620 45568
rect 22928 45620 22980 45626
rect 22928 45562 22980 45568
rect 24872 45558 24900 45834
rect 25332 45558 25360 46446
rect 18512 45552 18564 45558
rect 18512 45494 18564 45500
rect 24860 45552 24912 45558
rect 24860 45494 24912 45500
rect 25320 45552 25372 45558
rect 25320 45494 25372 45500
rect 15568 45484 15620 45490
rect 15568 45426 15620 45432
rect 14372 44940 14424 44946
rect 14372 44882 14424 44888
rect 15580 44538 15608 45426
rect 15568 44532 15620 44538
rect 15568 44474 15620 44480
rect 16948 41132 17000 41138
rect 16948 41074 17000 41080
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 16684 26382 16712 26930
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12544 17678 12572 25230
rect 16776 21418 16804 28154
rect 16960 27130 16988 41074
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17788 28490 17816 29106
rect 17132 28484 17184 28490
rect 17132 28426 17184 28432
rect 17776 28484 17828 28490
rect 17776 28426 17828 28432
rect 17144 28218 17172 28426
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17788 28082 17816 28426
rect 18156 28150 18184 33934
rect 18524 28626 18552 45494
rect 26252 45490 26280 46446
rect 27080 46442 27108 49200
rect 27620 47184 27672 47190
rect 27620 47126 27672 47132
rect 27068 46436 27120 46442
rect 27068 46378 27120 46384
rect 26976 45960 27028 45966
rect 26976 45902 27028 45908
rect 26988 45490 27016 45902
rect 27160 45892 27212 45898
rect 27160 45834 27212 45840
rect 22836 45484 22888 45490
rect 22836 45426 22888 45432
rect 24492 45484 24544 45490
rect 24492 45426 24544 45432
rect 26240 45484 26292 45490
rect 26240 45426 26292 45432
rect 26976 45484 27028 45490
rect 26976 45426 27028 45432
rect 22848 44810 22876 45426
rect 22836 44804 22888 44810
rect 22836 44746 22888 44752
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18512 28620 18564 28626
rect 18512 28562 18564 28568
rect 18788 28620 18840 28626
rect 18788 28562 18840 28568
rect 18144 28144 18196 28150
rect 18144 28086 18196 28092
rect 18420 28144 18472 28150
rect 18420 28086 18472 28092
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 17776 28076 17828 28082
rect 17776 28018 17828 28024
rect 17052 27470 17080 28018
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 17316 27396 17368 27402
rect 17316 27338 17368 27344
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 17052 26450 17080 27066
rect 17040 26444 17092 26450
rect 17040 26386 17092 26392
rect 17052 26234 17080 26386
rect 17328 26314 17356 27338
rect 18064 26994 18092 27406
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17868 26920 17920 26926
rect 17868 26862 17920 26868
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 16960 26206 17080 26234
rect 16960 23118 16988 26206
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 13648 17882 13676 18158
rect 15120 17882 15148 18158
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10428 3602 10456 3878
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9692 3126 9720 3470
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10704 3194 10732 3402
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 10980 800 11008 3538
rect 12360 3058 12388 4014
rect 12820 3738 12848 4014
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12912 800 12940 4014
rect 13096 2990 13124 17614
rect 17236 5710 17264 22102
rect 17328 19854 17356 26250
rect 17880 22778 17908 26862
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17880 22166 17908 22714
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14108 3738 14136 4762
rect 17328 4622 17356 19790
rect 18432 11762 18460 28086
rect 18604 27396 18656 27402
rect 18604 27338 18656 27344
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14108 3534 14136 3674
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13464 3058 13492 3470
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3126 13676 3334
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 17144 3058 17172 3878
rect 17880 3670 17908 5646
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 18616 3398 18644 27338
rect 18800 25362 18828 28562
rect 18788 25356 18840 25362
rect 18788 25298 18840 25304
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 17328 3126 17356 3334
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13556 800 13584 2858
rect 17420 800 17448 2926
rect 18800 2854 18828 25298
rect 18892 3194 18920 29242
rect 19996 28762 20024 36110
rect 20444 36032 20496 36038
rect 20444 35974 20496 35980
rect 19984 28756 20036 28762
rect 19984 28698 20036 28704
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10062 20024 28698
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 20076 9988 20128 9994
rect 20076 9930 20128 9936
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20088 4622 20116 9930
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19352 4078 19380 4422
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 18880 3188 18932 3194
rect 18880 3130 18932 3136
rect 19444 3074 19472 4014
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 3126 20024 4422
rect 20088 3602 20116 4558
rect 20456 4554 20484 35974
rect 22848 35894 22876 44746
rect 23848 40452 23900 40458
rect 23848 40394 23900 40400
rect 23480 40384 23532 40390
rect 23480 40326 23532 40332
rect 23492 40118 23520 40326
rect 23860 40186 23888 40394
rect 24400 40384 24452 40390
rect 24400 40326 24452 40332
rect 24504 40338 24532 45426
rect 26056 45348 26108 45354
rect 26056 45290 26108 45296
rect 25964 41064 26016 41070
rect 25964 41006 26016 41012
rect 24584 40996 24636 41002
rect 24584 40938 24636 40944
rect 24596 40526 24624 40938
rect 25320 40928 25372 40934
rect 25320 40870 25372 40876
rect 25332 40526 25360 40870
rect 25976 40730 26004 41006
rect 25964 40724 26016 40730
rect 25964 40666 26016 40672
rect 24584 40520 24636 40526
rect 24584 40462 24636 40468
rect 24860 40520 24912 40526
rect 24860 40462 24912 40468
rect 25320 40520 25372 40526
rect 25320 40462 25372 40468
rect 23848 40180 23900 40186
rect 23848 40122 23900 40128
rect 23480 40112 23532 40118
rect 23480 40054 23532 40060
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 23676 39370 23704 39782
rect 23664 39364 23716 39370
rect 23664 39306 23716 39312
rect 22848 35866 22968 35894
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22664 29102 22692 29582
rect 22652 29096 22704 29102
rect 22652 29038 22704 29044
rect 22664 28558 22692 29038
rect 22940 28966 22968 35866
rect 23860 31346 23888 40122
rect 24412 40118 24440 40326
rect 24504 40310 24624 40338
rect 24400 40112 24452 40118
rect 24400 40054 24452 40060
rect 24596 39098 24624 40310
rect 24872 39846 24900 40462
rect 24860 39840 24912 39846
rect 24860 39782 24912 39788
rect 24872 39370 24900 39782
rect 24860 39364 24912 39370
rect 24860 39306 24912 39312
rect 24584 39092 24636 39098
rect 24584 39034 24636 39040
rect 24308 36780 24360 36786
rect 24308 36722 24360 36728
rect 24320 35834 24348 36722
rect 24400 36576 24452 36582
rect 24400 36518 24452 36524
rect 24412 36174 24440 36518
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 24308 35828 24360 35834
rect 24308 35770 24360 35776
rect 24412 34610 24440 36110
rect 24400 34604 24452 34610
rect 24400 34546 24452 34552
rect 24492 34604 24544 34610
rect 24492 34546 24544 34552
rect 24412 33658 24440 34546
rect 24504 34202 24532 34546
rect 24492 34196 24544 34202
rect 24492 34138 24544 34144
rect 24400 33652 24452 33658
rect 24400 33594 24452 33600
rect 24412 31890 24440 33594
rect 24400 31884 24452 31890
rect 24400 31826 24452 31832
rect 24412 31346 24440 31826
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 24216 31340 24268 31346
rect 24216 31282 24268 31288
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 22928 28960 22980 28966
rect 22928 28902 22980 28908
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 22112 28082 22140 28358
rect 22848 28218 22876 28494
rect 22836 28212 22888 28218
rect 22836 28154 22888 28160
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 21916 27056 21968 27062
rect 21916 26998 21968 27004
rect 21928 24274 21956 26998
rect 22008 24744 22060 24750
rect 22008 24686 22060 24692
rect 21916 24268 21968 24274
rect 21916 24210 21968 24216
rect 22020 23866 22048 24686
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 22112 23186 22140 28018
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22572 26926 22600 27950
rect 22652 27872 22704 27878
rect 22652 27814 22704 27820
rect 22560 26920 22612 26926
rect 22560 26862 22612 26868
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22480 25294 22508 25638
rect 22664 25294 22692 27814
rect 23020 26920 23072 26926
rect 23020 26862 23072 26868
rect 23032 26382 23060 26862
rect 23216 26450 23244 29106
rect 23480 29028 23532 29034
rect 23480 28970 23532 28976
rect 23492 28082 23520 28970
rect 23756 28484 23808 28490
rect 23756 28426 23808 28432
rect 23768 28082 23796 28426
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23768 27606 23796 28018
rect 23756 27600 23808 27606
rect 23756 27542 23808 27548
rect 24122 27432 24178 27441
rect 24122 27367 24124 27376
rect 24176 27367 24178 27376
rect 24124 27338 24176 27344
rect 23204 26444 23256 26450
rect 23204 26386 23256 26392
rect 23020 26376 23072 26382
rect 23020 26318 23072 26324
rect 23216 25838 23244 26386
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 23492 25294 23520 25842
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 22744 25152 22796 25158
rect 22744 25094 22796 25100
rect 22928 25152 22980 25158
rect 22928 25094 22980 25100
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22204 24410 22232 24686
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22756 24138 22784 25094
rect 22940 24206 22968 25094
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 22744 24132 22796 24138
rect 22744 24074 22796 24080
rect 23124 24070 23152 25230
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 23308 24410 23336 25094
rect 23492 24818 23520 25230
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23296 24404 23348 24410
rect 23296 24346 23348 24352
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 23952 23662 23980 24142
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 23952 22710 23980 23598
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24136 20874 24164 21286
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 22112 4146 22140 10406
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21376 3194 21404 3402
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 19352 3046 19472 3074
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 22020 3058 22048 3470
rect 22008 3052 22060 3058
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 19352 800 19380 3046
rect 22008 2994 22060 3000
rect 22204 2990 22232 3878
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 19444 2650 19472 2926
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20640 800 20668 2926
rect 22572 800 22600 2926
rect 24228 2514 24256 31282
rect 24400 29504 24452 29510
rect 24400 29446 24452 29452
rect 24412 29170 24440 29446
rect 24596 29306 24624 39034
rect 24872 37806 24900 39306
rect 25688 39296 25740 39302
rect 25688 39238 25740 39244
rect 25596 38208 25648 38214
rect 25596 38150 25648 38156
rect 25608 37874 25636 38150
rect 25596 37868 25648 37874
rect 25596 37810 25648 37816
rect 24860 37800 24912 37806
rect 24860 37742 24912 37748
rect 24872 37312 24900 37742
rect 24780 37284 24900 37312
rect 24676 37120 24728 37126
rect 24676 37062 24728 37068
rect 24688 36174 24716 37062
rect 24780 36582 24808 37284
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 24768 36576 24820 36582
rect 24768 36518 24820 36524
rect 24676 36168 24728 36174
rect 24676 36110 24728 36116
rect 24964 35834 24992 37198
rect 25412 36576 25464 36582
rect 25412 36518 25464 36524
rect 24952 35828 25004 35834
rect 24952 35770 25004 35776
rect 24952 35692 25004 35698
rect 24952 35634 25004 35640
rect 25044 35692 25096 35698
rect 25044 35634 25096 35640
rect 24964 35290 24992 35634
rect 24952 35284 25004 35290
rect 24952 35226 25004 35232
rect 25056 35086 25084 35634
rect 25424 35630 25452 36518
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 25504 35624 25556 35630
rect 25504 35566 25556 35572
rect 25516 35086 25544 35566
rect 25700 35494 25728 39238
rect 26068 38554 26096 45290
rect 27172 45082 27200 45834
rect 27436 45416 27488 45422
rect 27436 45358 27488 45364
rect 27448 45082 27476 45358
rect 27160 45076 27212 45082
rect 27160 45018 27212 45024
rect 27436 45076 27488 45082
rect 27436 45018 27488 45024
rect 26700 44872 26752 44878
rect 26700 44814 26752 44820
rect 26608 41064 26660 41070
rect 26608 41006 26660 41012
rect 26620 39642 26648 41006
rect 26608 39636 26660 39642
rect 26608 39578 26660 39584
rect 26056 38548 26108 38554
rect 26056 38490 26108 38496
rect 25780 38344 25832 38350
rect 25780 38286 25832 38292
rect 25792 37466 25820 38286
rect 25780 37460 25832 37466
rect 25780 37402 25832 37408
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 25792 36378 25820 37198
rect 25780 36372 25832 36378
rect 25780 36314 25832 36320
rect 26712 36106 26740 44814
rect 27632 42702 27660 47126
rect 28000 47054 28028 49286
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 33478 49200 33590 50000
rect 34122 49200 34234 50000
rect 35410 49200 35522 50000
rect 36054 49200 36166 50000
rect 36698 49200 36810 50000
rect 37986 49200 38098 50000
rect 38630 49200 38742 50000
rect 39918 49200 40030 50000
rect 40562 49200 40674 50000
rect 41850 49314 41962 50000
rect 41850 49286 42104 49314
rect 41850 49200 41962 49286
rect 29656 47138 29684 49200
rect 28816 47116 28868 47122
rect 29656 47110 30236 47138
rect 28816 47058 28868 47064
rect 27988 47048 28040 47054
rect 27988 46990 28040 46996
rect 28828 45966 28856 47058
rect 29736 47048 29788 47054
rect 29736 46990 29788 46996
rect 29748 46578 29776 46990
rect 29736 46572 29788 46578
rect 29736 46514 29788 46520
rect 29920 46504 29972 46510
rect 29920 46446 29972 46452
rect 28816 45960 28868 45966
rect 28816 45902 28868 45908
rect 29736 45960 29788 45966
rect 29736 45902 29788 45908
rect 29748 45558 29776 45902
rect 29736 45552 29788 45558
rect 29736 45494 29788 45500
rect 29932 45082 29960 46446
rect 30208 45554 30236 47110
rect 30300 46510 30328 49200
rect 32772 47048 32824 47054
rect 32772 46990 32824 46996
rect 32784 46578 32812 46990
rect 32772 46572 32824 46578
rect 32772 46514 32824 46520
rect 33520 46510 33548 49200
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 35808 46572 35860 46578
rect 35808 46514 35860 46520
rect 30288 46504 30340 46510
rect 30288 46446 30340 46452
rect 32956 46504 33008 46510
rect 32956 46446 33008 46452
rect 33508 46504 33560 46510
rect 33508 46446 33560 46452
rect 32968 46170 32996 46446
rect 35716 46436 35768 46442
rect 35716 46378 35768 46384
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 32956 46164 33008 46170
rect 32956 46106 33008 46112
rect 35728 45966 35756 46378
rect 32772 45960 32824 45966
rect 32772 45902 32824 45908
rect 35716 45960 35768 45966
rect 35716 45902 35768 45908
rect 32784 45626 32812 45902
rect 35820 45830 35848 46514
rect 35900 46368 35952 46374
rect 35900 46310 35952 46316
rect 35912 45898 35940 46310
rect 36096 46034 36124 49200
rect 36740 46442 36768 49200
rect 38672 47462 38700 49200
rect 38660 47456 38712 47462
rect 38660 47398 38712 47404
rect 39948 47456 40000 47462
rect 39948 47398 40000 47404
rect 37280 47048 37332 47054
rect 37280 46990 37332 46996
rect 37292 46578 37320 46990
rect 37280 46572 37332 46578
rect 37280 46514 37332 46520
rect 37464 46504 37516 46510
rect 37464 46446 37516 46452
rect 36728 46436 36780 46442
rect 36728 46378 36780 46384
rect 36084 46028 36136 46034
rect 36084 45970 36136 45976
rect 35900 45892 35952 45898
rect 35900 45834 35952 45840
rect 35808 45824 35860 45830
rect 35808 45766 35860 45772
rect 32772 45620 32824 45626
rect 32772 45562 32824 45568
rect 30208 45526 30328 45554
rect 30300 45422 30328 45526
rect 30288 45416 30340 45422
rect 30288 45358 30340 45364
rect 29920 45076 29972 45082
rect 29920 45018 29972 45024
rect 29920 44872 29972 44878
rect 29920 44814 29972 44820
rect 29932 44470 29960 44814
rect 29920 44464 29972 44470
rect 29920 44406 29972 44412
rect 32784 44334 32812 45562
rect 36084 45484 36136 45490
rect 36084 45426 36136 45432
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 32772 44328 32824 44334
rect 32772 44270 32824 44276
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 30656 42764 30708 42770
rect 30656 42706 30708 42712
rect 27620 42696 27672 42702
rect 27620 42638 27672 42644
rect 27160 42560 27212 42566
rect 27160 42502 27212 42508
rect 28540 42560 28592 42566
rect 28540 42502 28592 42508
rect 27172 42226 27200 42502
rect 28552 42226 28580 42502
rect 27160 42220 27212 42226
rect 27160 42162 27212 42168
rect 28540 42220 28592 42226
rect 28540 42162 28592 42168
rect 26976 42016 27028 42022
rect 26976 41958 27028 41964
rect 29644 42016 29696 42022
rect 29644 41958 29696 41964
rect 26988 41546 27016 41958
rect 29656 41614 29684 41958
rect 29552 41608 29604 41614
rect 29552 41550 29604 41556
rect 29644 41608 29696 41614
rect 29644 41550 29696 41556
rect 26976 41540 27028 41546
rect 26976 41482 27028 41488
rect 27896 41472 27948 41478
rect 27896 41414 27948 41420
rect 27068 41132 27120 41138
rect 27068 41074 27120 41080
rect 27080 40526 27108 41074
rect 27908 40730 27936 41414
rect 29000 41132 29052 41138
rect 29000 41074 29052 41080
rect 29012 40730 29040 41074
rect 29368 40928 29420 40934
rect 29368 40870 29420 40876
rect 27896 40724 27948 40730
rect 27816 40684 27896 40712
rect 27252 40656 27304 40662
rect 27252 40598 27304 40604
rect 27068 40520 27120 40526
rect 27068 40462 27120 40468
rect 27080 39642 27108 40462
rect 27264 40118 27292 40598
rect 27712 40452 27764 40458
rect 27712 40394 27764 40400
rect 27252 40112 27304 40118
rect 27252 40054 27304 40060
rect 27068 39636 27120 39642
rect 27068 39578 27120 39584
rect 27080 39438 27108 39578
rect 27068 39432 27120 39438
rect 27068 39374 27120 39380
rect 27080 39114 27108 39374
rect 27724 39370 27752 40394
rect 27712 39364 27764 39370
rect 27712 39306 27764 39312
rect 27816 39302 27844 40684
rect 27896 40666 27948 40672
rect 29000 40724 29052 40730
rect 29000 40666 29052 40672
rect 29380 40526 29408 40870
rect 29564 40594 29592 41550
rect 30012 41132 30064 41138
rect 30012 41074 30064 41080
rect 29552 40588 29604 40594
rect 29552 40530 29604 40536
rect 27896 40520 27948 40526
rect 27896 40462 27948 40468
rect 27988 40520 28040 40526
rect 27988 40462 28040 40468
rect 29368 40520 29420 40526
rect 29368 40462 29420 40468
rect 27908 39846 27936 40462
rect 28000 40186 28028 40462
rect 29184 40452 29236 40458
rect 29184 40394 29236 40400
rect 28172 40384 28224 40390
rect 28172 40326 28224 40332
rect 27988 40180 28040 40186
rect 27988 40122 28040 40128
rect 27896 39840 27948 39846
rect 27896 39782 27948 39788
rect 27908 39438 27936 39782
rect 28000 39574 28028 40122
rect 27988 39568 28040 39574
rect 27988 39510 28040 39516
rect 27896 39432 27948 39438
rect 27896 39374 27948 39380
rect 27804 39296 27856 39302
rect 27804 39238 27856 39244
rect 26988 39086 27108 39114
rect 26792 37664 26844 37670
rect 26792 37606 26844 37612
rect 26804 37330 26832 37606
rect 26792 37324 26844 37330
rect 26792 37266 26844 37272
rect 26988 37262 27016 39086
rect 28184 38350 28212 40326
rect 29196 40050 29224 40394
rect 29564 40118 29592 40530
rect 30024 40458 30052 41074
rect 30012 40452 30064 40458
rect 30012 40394 30064 40400
rect 29552 40112 29604 40118
rect 29552 40054 29604 40060
rect 29184 40044 29236 40050
rect 29184 39986 29236 39992
rect 30024 39846 30052 40394
rect 30196 40044 30248 40050
rect 30196 39986 30248 39992
rect 30012 39840 30064 39846
rect 30012 39782 30064 39788
rect 28540 39296 28592 39302
rect 28540 39238 28592 39244
rect 28172 38344 28224 38350
rect 28172 38286 28224 38292
rect 27620 37936 27672 37942
rect 27620 37878 27672 37884
rect 27068 37324 27120 37330
rect 27068 37266 27120 37272
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 27080 36666 27108 37266
rect 27252 37120 27304 37126
rect 27252 37062 27304 37068
rect 27264 36786 27292 37062
rect 27632 36854 27660 37878
rect 28552 37262 28580 39238
rect 30024 38962 30052 39782
rect 30208 39438 30236 39986
rect 30196 39432 30248 39438
rect 30196 39374 30248 39380
rect 30012 38956 30064 38962
rect 30012 38898 30064 38904
rect 30196 38888 30248 38894
rect 30196 38830 30248 38836
rect 29828 38752 29880 38758
rect 29828 38694 29880 38700
rect 29552 38412 29604 38418
rect 29552 38354 29604 38360
rect 28908 38208 28960 38214
rect 28908 38150 28960 38156
rect 28920 37262 28948 38150
rect 29460 37868 29512 37874
rect 29460 37810 29512 37816
rect 29472 37466 29500 37810
rect 29460 37460 29512 37466
rect 29460 37402 29512 37408
rect 29564 37398 29592 38354
rect 29736 38276 29788 38282
rect 29736 38218 29788 38224
rect 29748 37874 29776 38218
rect 29736 37868 29788 37874
rect 29736 37810 29788 37816
rect 29552 37392 29604 37398
rect 29552 37334 29604 37340
rect 29000 37324 29052 37330
rect 29000 37266 29052 37272
rect 28540 37256 28592 37262
rect 28540 37198 28592 37204
rect 28908 37256 28960 37262
rect 28908 37198 28960 37204
rect 28724 37188 28776 37194
rect 28724 37130 28776 37136
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 28368 36854 28396 37062
rect 27620 36848 27672 36854
rect 27620 36790 27672 36796
rect 27896 36848 27948 36854
rect 27896 36790 27948 36796
rect 28356 36848 28408 36854
rect 28356 36790 28408 36796
rect 27252 36780 27304 36786
rect 27252 36722 27304 36728
rect 27080 36638 27384 36666
rect 26884 36372 26936 36378
rect 26884 36314 26936 36320
rect 26792 36168 26844 36174
rect 26792 36110 26844 36116
rect 26700 36100 26752 36106
rect 26700 36042 26752 36048
rect 26056 35760 26108 35766
rect 26056 35702 26108 35708
rect 25872 35692 25924 35698
rect 25872 35634 25924 35640
rect 25688 35488 25740 35494
rect 25688 35430 25740 35436
rect 25044 35080 25096 35086
rect 25044 35022 25096 35028
rect 25504 35080 25556 35086
rect 25504 35022 25556 35028
rect 24860 35012 24912 35018
rect 24860 34954 24912 34960
rect 24872 33998 24900 34954
rect 25412 34740 25464 34746
rect 25412 34682 25464 34688
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 24872 32978 24900 33934
rect 24860 32972 24912 32978
rect 24860 32914 24912 32920
rect 25424 32910 25452 34682
rect 25516 33658 25544 35022
rect 25884 35018 25912 35634
rect 25964 35488 26016 35494
rect 25964 35430 26016 35436
rect 25872 35012 25924 35018
rect 25872 34954 25924 34960
rect 25884 34746 25912 34954
rect 25976 34950 26004 35430
rect 26068 35154 26096 35702
rect 26804 35562 26832 36110
rect 26896 36038 26924 36314
rect 26884 36032 26936 36038
rect 26884 35974 26936 35980
rect 27080 35766 27108 36638
rect 27160 36576 27212 36582
rect 27160 36518 27212 36524
rect 27172 36174 27200 36518
rect 27252 36304 27304 36310
rect 27252 36246 27304 36252
rect 27160 36168 27212 36174
rect 27160 36110 27212 36116
rect 27068 35760 27120 35766
rect 27068 35702 27120 35708
rect 27172 35630 27200 36110
rect 27264 35698 27292 36246
rect 27356 36174 27384 36638
rect 27344 36168 27396 36174
rect 27344 36110 27396 36116
rect 27804 36032 27856 36038
rect 27804 35974 27856 35980
rect 27252 35692 27304 35698
rect 27252 35634 27304 35640
rect 27160 35624 27212 35630
rect 27160 35566 27212 35572
rect 26792 35556 26844 35562
rect 26792 35498 26844 35504
rect 26148 35488 26200 35494
rect 26148 35430 26200 35436
rect 27068 35488 27120 35494
rect 27068 35430 27120 35436
rect 26056 35148 26108 35154
rect 26056 35090 26108 35096
rect 25964 34944 26016 34950
rect 25964 34886 26016 34892
rect 25872 34740 25924 34746
rect 25872 34682 25924 34688
rect 25976 33930 26004 34886
rect 25964 33924 26016 33930
rect 25964 33866 26016 33872
rect 25504 33652 25556 33658
rect 25504 33594 25556 33600
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 26068 32842 26096 35090
rect 26160 34746 26188 35430
rect 26148 34740 26200 34746
rect 26148 34682 26200 34688
rect 27080 34610 27108 35430
rect 27816 35086 27844 35974
rect 27804 35080 27856 35086
rect 27804 35022 27856 35028
rect 27528 34944 27580 34950
rect 27528 34886 27580 34892
rect 27540 34678 27568 34886
rect 27528 34672 27580 34678
rect 27528 34614 27580 34620
rect 27908 34610 27936 36790
rect 28736 35562 28764 37130
rect 28724 35556 28776 35562
rect 28724 35498 28776 35504
rect 27988 35012 28040 35018
rect 27988 34954 28040 34960
rect 28000 34746 28028 34954
rect 28736 34950 28764 35498
rect 29012 35494 29040 37266
rect 29840 37262 29868 38694
rect 30208 38214 30236 38830
rect 30104 38208 30156 38214
rect 30104 38150 30156 38156
rect 30196 38208 30248 38214
rect 30196 38150 30248 38156
rect 30116 38010 30144 38150
rect 30104 38004 30156 38010
rect 30104 37946 30156 37952
rect 30208 37942 30236 38150
rect 30196 37936 30248 37942
rect 30196 37878 30248 37884
rect 29828 37256 29880 37262
rect 29828 37198 29880 37204
rect 30196 36576 30248 36582
rect 30196 36518 30248 36524
rect 30208 36242 30236 36518
rect 29184 36236 29236 36242
rect 29184 36178 29236 36184
rect 30196 36236 30248 36242
rect 30196 36178 30248 36184
rect 29000 35488 29052 35494
rect 29000 35430 29052 35436
rect 29000 35080 29052 35086
rect 29000 35022 29052 35028
rect 28724 34944 28776 34950
rect 28724 34886 28776 34892
rect 27988 34740 28040 34746
rect 27988 34682 28040 34688
rect 27068 34604 27120 34610
rect 27068 34546 27120 34552
rect 27896 34604 27948 34610
rect 27896 34546 27948 34552
rect 27908 34202 27936 34546
rect 27620 34196 27672 34202
rect 27620 34138 27672 34144
rect 27896 34196 27948 34202
rect 27896 34138 27948 34144
rect 26148 33516 26200 33522
rect 26148 33458 26200 33464
rect 26160 33114 26188 33458
rect 26148 33108 26200 33114
rect 26148 33050 26200 33056
rect 27632 32978 27660 34138
rect 28632 33924 28684 33930
rect 28632 33866 28684 33872
rect 28644 33522 28672 33866
rect 29012 33862 29040 35022
rect 29000 33856 29052 33862
rect 29000 33798 29052 33804
rect 28632 33516 28684 33522
rect 28632 33458 28684 33464
rect 27620 32972 27672 32978
rect 27620 32914 27672 32920
rect 29012 32910 29040 33798
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 26056 32836 26108 32842
rect 26056 32778 26108 32784
rect 25320 32768 25372 32774
rect 25320 32710 25372 32716
rect 25332 32434 25360 32710
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 24952 32224 25004 32230
rect 24952 32166 25004 32172
rect 24964 31822 24992 32166
rect 26068 32026 26096 32778
rect 28816 32768 28868 32774
rect 28816 32710 28868 32716
rect 28828 32502 28856 32710
rect 28816 32496 28868 32502
rect 28816 32438 28868 32444
rect 29196 32450 29224 36178
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 29564 35698 29592 35974
rect 30668 35894 30696 42706
rect 33784 42696 33836 42702
rect 33784 42638 33836 42644
rect 33508 42560 33560 42566
rect 33508 42502 33560 42508
rect 33520 42294 33548 42502
rect 33508 42288 33560 42294
rect 33508 42230 33560 42236
rect 31392 42220 31444 42226
rect 31392 42162 31444 42168
rect 32680 42220 32732 42226
rect 32680 42162 32732 42168
rect 31208 42016 31260 42022
rect 31208 41958 31260 41964
rect 31220 41546 31248 41958
rect 31208 41540 31260 41546
rect 31208 41482 31260 41488
rect 30932 41472 30984 41478
rect 30932 41414 30984 41420
rect 30944 41070 30972 41414
rect 31404 41274 31432 42162
rect 32496 42016 32548 42022
rect 32496 41958 32548 41964
rect 31392 41268 31444 41274
rect 31392 41210 31444 41216
rect 32508 41206 32536 41958
rect 32692 41818 32720 42162
rect 33140 42152 33192 42158
rect 33140 42094 33192 42100
rect 32680 41812 32732 41818
rect 32680 41754 32732 41760
rect 33152 41614 33180 42094
rect 33140 41608 33192 41614
rect 33140 41550 33192 41556
rect 33600 41608 33652 41614
rect 33600 41550 33652 41556
rect 32496 41200 32548 41206
rect 32496 41142 32548 41148
rect 30932 41064 30984 41070
rect 30932 41006 30984 41012
rect 33152 40934 33180 41550
rect 33140 40928 33192 40934
rect 33140 40870 33192 40876
rect 32588 40724 32640 40730
rect 32588 40666 32640 40672
rect 30748 40384 30800 40390
rect 30748 40326 30800 40332
rect 30760 39438 30788 40326
rect 31760 40044 31812 40050
rect 31760 39986 31812 39992
rect 31024 39908 31076 39914
rect 31024 39850 31076 39856
rect 30748 39432 30800 39438
rect 30748 39374 30800 39380
rect 30840 39432 30892 39438
rect 30840 39374 30892 39380
rect 30760 38350 30788 39374
rect 30852 39030 30880 39374
rect 31036 39098 31064 39850
rect 31772 39438 31800 39986
rect 32600 39642 32628 40666
rect 33612 40526 33640 41550
rect 33692 40928 33744 40934
rect 33692 40870 33744 40876
rect 33600 40520 33652 40526
rect 33600 40462 33652 40468
rect 32588 39636 32640 39642
rect 32588 39578 32640 39584
rect 31760 39432 31812 39438
rect 31760 39374 31812 39380
rect 31484 39296 31536 39302
rect 31484 39238 31536 39244
rect 31024 39092 31076 39098
rect 31024 39034 31076 39040
rect 30840 39024 30892 39030
rect 30840 38966 30892 38972
rect 30932 38888 30984 38894
rect 30932 38830 30984 38836
rect 30748 38344 30800 38350
rect 30748 38286 30800 38292
rect 30760 37670 30788 38286
rect 30748 37664 30800 37670
rect 30748 37606 30800 37612
rect 30944 37194 30972 38830
rect 31496 38282 31524 39238
rect 31772 38894 31800 39374
rect 31852 39024 31904 39030
rect 31852 38966 31904 38972
rect 31760 38888 31812 38894
rect 31760 38830 31812 38836
rect 31484 38276 31536 38282
rect 31484 38218 31536 38224
rect 31300 38208 31352 38214
rect 31300 38150 31352 38156
rect 31312 37874 31340 38150
rect 31300 37868 31352 37874
rect 31300 37810 31352 37816
rect 31864 37194 31892 38966
rect 33704 38894 33732 40870
rect 33796 40730 33824 42638
rect 34520 42016 34572 42022
rect 34520 41958 34572 41964
rect 35348 42016 35400 42022
rect 35348 41958 35400 41964
rect 35808 42016 35860 42022
rect 35808 41958 35860 41964
rect 34428 41268 34480 41274
rect 34428 41210 34480 41216
rect 33874 41032 33930 41041
rect 34440 41002 34468 41210
rect 34532 41206 34560 41958
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34612 41540 34664 41546
rect 34612 41482 34664 41488
rect 34520 41200 34572 41206
rect 34520 41142 34572 41148
rect 34624 41188 34652 41482
rect 34704 41200 34756 41206
rect 34624 41160 34704 41188
rect 33874 40967 33876 40976
rect 33928 40967 33930 40976
rect 34428 40996 34480 41002
rect 33876 40938 33928 40944
rect 34428 40938 34480 40944
rect 33784 40724 33836 40730
rect 33784 40666 33836 40672
rect 33888 40458 33916 40938
rect 34624 40934 34652 41160
rect 34704 41142 34756 41148
rect 34796 41132 34848 41138
rect 34796 41074 34848 41080
rect 34808 41041 34836 41074
rect 35360 41070 35388 41958
rect 35820 41614 35848 41958
rect 35808 41608 35860 41614
rect 35808 41550 35860 41556
rect 35348 41064 35400 41070
rect 34794 41032 34850 41041
rect 35348 41006 35400 41012
rect 34794 40967 34850 40976
rect 34612 40928 34664 40934
rect 34612 40870 34664 40876
rect 34796 40928 34848 40934
rect 34796 40870 34848 40876
rect 35716 40928 35768 40934
rect 35716 40870 35768 40876
rect 33876 40452 33928 40458
rect 33876 40394 33928 40400
rect 34808 39438 34836 40870
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35728 40526 35756 40870
rect 35716 40520 35768 40526
rect 35716 40462 35768 40468
rect 35348 40384 35400 40390
rect 35348 40326 35400 40332
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35360 39438 35388 40326
rect 35900 40180 35952 40186
rect 35900 40122 35952 40128
rect 35912 39506 35940 40122
rect 35900 39500 35952 39506
rect 35900 39442 35952 39448
rect 34796 39432 34848 39438
rect 34796 39374 34848 39380
rect 35348 39432 35400 39438
rect 35348 39374 35400 39380
rect 35440 39432 35492 39438
rect 35440 39374 35492 39380
rect 34796 39296 34848 39302
rect 34796 39238 34848 39244
rect 32220 38888 32272 38894
rect 32220 38830 32272 38836
rect 33692 38888 33744 38894
rect 33692 38830 33744 38836
rect 32232 38486 32260 38830
rect 32864 38752 32916 38758
rect 32864 38694 32916 38700
rect 32220 38480 32272 38486
rect 32220 38422 32272 38428
rect 32128 38344 32180 38350
rect 32128 38286 32180 38292
rect 32140 37806 32168 38286
rect 32232 38214 32260 38422
rect 32876 38350 32904 38694
rect 33704 38418 33732 38830
rect 33692 38412 33744 38418
rect 33692 38354 33744 38360
rect 34808 38350 34836 39238
rect 35452 39098 35480 39374
rect 35440 39092 35492 39098
rect 35440 39034 35492 39040
rect 35348 38888 35400 38894
rect 35348 38830 35400 38836
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 32864 38344 32916 38350
rect 32864 38286 32916 38292
rect 34796 38344 34848 38350
rect 34796 38286 34848 38292
rect 35360 38214 35388 38830
rect 35624 38752 35676 38758
rect 35624 38694 35676 38700
rect 32220 38208 32272 38214
rect 32220 38150 32272 38156
rect 32680 38208 32732 38214
rect 32680 38150 32732 38156
rect 35348 38208 35400 38214
rect 35348 38150 35400 38156
rect 32692 37942 32720 38150
rect 32680 37936 32732 37942
rect 32680 37878 32732 37884
rect 35360 37806 35388 38150
rect 35636 38010 35664 38694
rect 35624 38004 35676 38010
rect 35624 37946 35676 37952
rect 35636 37806 35664 37946
rect 35716 37868 35768 37874
rect 35716 37810 35768 37816
rect 32128 37800 32180 37806
rect 32128 37742 32180 37748
rect 35348 37800 35400 37806
rect 35348 37742 35400 37748
rect 35624 37800 35676 37806
rect 35624 37742 35676 37748
rect 30932 37188 30984 37194
rect 30932 37130 30984 37136
rect 31852 37188 31904 37194
rect 31852 37130 31904 37136
rect 30944 36174 30972 37130
rect 32140 36718 32168 37742
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35360 37330 35388 37742
rect 35636 37398 35664 37742
rect 35624 37392 35676 37398
rect 35624 37334 35676 37340
rect 35348 37324 35400 37330
rect 35348 37266 35400 37272
rect 35728 37262 35756 37810
rect 35992 37664 36044 37670
rect 35992 37606 36044 37612
rect 35716 37256 35768 37262
rect 35716 37198 35768 37204
rect 35440 37120 35492 37126
rect 35440 37062 35492 37068
rect 33140 36780 33192 36786
rect 33140 36722 33192 36728
rect 31760 36712 31812 36718
rect 31760 36654 31812 36660
rect 32128 36712 32180 36718
rect 32128 36654 32180 36660
rect 30932 36168 30984 36174
rect 30932 36110 30984 36116
rect 30668 35866 30880 35894
rect 29552 35692 29604 35698
rect 29552 35634 29604 35640
rect 29368 35488 29420 35494
rect 29368 35430 29420 35436
rect 29380 34678 29408 35430
rect 29368 34672 29420 34678
rect 29368 34614 29420 34620
rect 29736 34536 29788 34542
rect 29736 34478 29788 34484
rect 29276 34400 29328 34406
rect 29276 34342 29328 34348
rect 29288 32978 29316 34342
rect 29748 33454 29776 34478
rect 30380 33992 30432 33998
rect 30380 33934 30432 33940
rect 30656 33992 30708 33998
rect 30656 33934 30708 33940
rect 29736 33448 29788 33454
rect 29736 33390 29788 33396
rect 30392 33114 30420 33934
rect 30668 33114 30696 33934
rect 30380 33108 30432 33114
rect 30380 33050 30432 33056
rect 30656 33108 30708 33114
rect 30656 33050 30708 33056
rect 29276 32972 29328 32978
rect 29276 32914 29328 32920
rect 29552 32972 29604 32978
rect 29552 32914 29604 32920
rect 29564 32570 29592 32914
rect 30380 32836 30432 32842
rect 30380 32778 30432 32784
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29736 32564 29788 32570
rect 29736 32506 29788 32512
rect 28828 32366 28856 32438
rect 29196 32434 29316 32450
rect 29184 32428 29316 32434
rect 29236 32422 29316 32428
rect 29184 32370 29236 32376
rect 27620 32360 27672 32366
rect 27620 32302 27672 32308
rect 28816 32360 28868 32366
rect 28816 32302 28868 32308
rect 26056 32020 26108 32026
rect 26056 31962 26108 31968
rect 27632 31890 27660 32302
rect 27804 32292 27856 32298
rect 27804 32234 27856 32240
rect 29184 32292 29236 32298
rect 29184 32234 29236 32240
rect 27620 31884 27672 31890
rect 27620 31826 27672 31832
rect 27816 31822 27844 32234
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 24952 31816 25004 31822
rect 24952 31758 25004 31764
rect 27804 31816 27856 31822
rect 27804 31758 27856 31764
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 27988 31680 28040 31686
rect 27988 31622 28040 31628
rect 25136 31340 25188 31346
rect 25136 31282 25188 31288
rect 24860 31136 24912 31142
rect 24860 31078 24912 31084
rect 24872 30734 24900 31078
rect 25148 30938 25176 31282
rect 28000 31210 28028 31622
rect 27988 31204 28040 31210
rect 27988 31146 28040 31152
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 27436 30592 27488 30598
rect 27436 30534 27488 30540
rect 24676 29640 24728 29646
rect 24676 29582 24728 29588
rect 24860 29640 24912 29646
rect 25596 29640 25648 29646
rect 24912 29600 24992 29628
rect 24860 29582 24912 29588
rect 24688 29306 24716 29582
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24860 29504 24912 29510
rect 24860 29446 24912 29452
rect 24584 29300 24636 29306
rect 24584 29242 24636 29248
rect 24676 29300 24728 29306
rect 24676 29242 24728 29248
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 24780 28694 24808 29446
rect 24872 29238 24900 29446
rect 24860 29232 24912 29238
rect 24860 29174 24912 29180
rect 24768 28688 24820 28694
rect 24768 28630 24820 28636
rect 24872 25838 24900 29174
rect 24964 28762 24992 29600
rect 25594 29608 25596 29617
rect 26332 29640 26384 29646
rect 25648 29608 25650 29617
rect 26332 29582 26384 29588
rect 25594 29543 25650 29552
rect 25872 29572 25924 29578
rect 25872 29514 25924 29520
rect 25884 29306 25912 29514
rect 25964 29504 26016 29510
rect 25964 29446 26016 29452
rect 25872 29300 25924 29306
rect 25872 29242 25924 29248
rect 25872 29164 25924 29170
rect 25976 29152 26004 29446
rect 26240 29300 26292 29306
rect 26240 29242 26292 29248
rect 25924 29124 26004 29152
rect 25872 29106 25924 29112
rect 25780 29096 25832 29102
rect 25778 29064 25780 29073
rect 25832 29064 25834 29073
rect 25778 28999 25834 29008
rect 24952 28756 25004 28762
rect 24952 28698 25004 28704
rect 25320 28552 25372 28558
rect 25320 28494 25372 28500
rect 25228 27940 25280 27946
rect 25228 27882 25280 27888
rect 24952 27872 25004 27878
rect 24952 27814 25004 27820
rect 24964 26926 24992 27814
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25148 26994 25176 27406
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 25136 26852 25188 26858
rect 25136 26794 25188 26800
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 24780 24070 24808 24754
rect 24872 24138 24900 25774
rect 25148 25294 25176 26794
rect 25240 26450 25268 27882
rect 25228 26444 25280 26450
rect 25228 26386 25280 26392
rect 25332 25294 25360 28494
rect 25976 28014 26004 29124
rect 26146 29064 26202 29073
rect 26056 29028 26108 29034
rect 26146 28999 26202 29008
rect 26056 28970 26108 28976
rect 26068 28558 26096 28970
rect 26160 28762 26188 28999
rect 26252 28762 26280 29242
rect 26344 29170 26372 29582
rect 27448 29170 27476 30534
rect 28078 29608 28134 29617
rect 28078 29543 28134 29552
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 26332 29164 26384 29170
rect 26332 29106 26384 29112
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 26700 28960 26752 28966
rect 26700 28902 26752 28908
rect 26712 28762 26740 28902
rect 26148 28756 26200 28762
rect 26148 28698 26200 28704
rect 26240 28756 26292 28762
rect 26240 28698 26292 28704
rect 26700 28756 26752 28762
rect 26700 28698 26752 28704
rect 26148 28620 26200 28626
rect 26148 28562 26200 28568
rect 26056 28552 26108 28558
rect 26056 28494 26108 28500
rect 26160 28082 26188 28562
rect 27448 28558 27476 29106
rect 27632 29050 27660 29242
rect 28092 29170 28120 29543
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 27540 29022 27660 29050
rect 27540 28966 27568 29022
rect 27528 28960 27580 28966
rect 27528 28902 27580 28908
rect 28184 28762 28212 29106
rect 28172 28756 28224 28762
rect 28172 28698 28224 28704
rect 26332 28552 26384 28558
rect 26332 28494 26384 28500
rect 27436 28552 27488 28558
rect 27436 28494 27488 28500
rect 26344 28218 26372 28494
rect 27448 28218 27476 28494
rect 27620 28416 27672 28422
rect 27620 28358 27672 28364
rect 26332 28212 26384 28218
rect 26332 28154 26384 28160
rect 27436 28212 27488 28218
rect 27436 28154 27488 28160
rect 26148 28076 26200 28082
rect 26148 28018 26200 28024
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 25964 28008 26016 28014
rect 25964 27950 26016 27956
rect 25504 27532 25556 27538
rect 25504 27474 25556 27480
rect 25516 27334 25544 27474
rect 25596 27464 25648 27470
rect 25596 27406 25648 27412
rect 25504 27328 25556 27334
rect 25504 27270 25556 27276
rect 25412 27056 25464 27062
rect 25412 26998 25464 27004
rect 25424 26586 25452 26998
rect 25608 26586 25636 27406
rect 25780 26920 25832 26926
rect 25780 26862 25832 26868
rect 25412 26580 25464 26586
rect 25412 26522 25464 26528
rect 25596 26580 25648 26586
rect 25596 26522 25648 26528
rect 25792 26382 25820 26862
rect 25976 26586 26004 27950
rect 26160 27674 26188 28018
rect 26148 27668 26200 27674
rect 26148 27610 26200 27616
rect 26436 27606 26464 28018
rect 26056 27600 26108 27606
rect 26056 27542 26108 27548
rect 26424 27600 26476 27606
rect 26424 27542 26476 27548
rect 26516 27600 26568 27606
rect 26516 27542 26568 27548
rect 26068 27470 26096 27542
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 26436 26858 26464 27542
rect 26528 27441 26556 27542
rect 27172 27470 27200 28018
rect 27160 27464 27212 27470
rect 26514 27432 26570 27441
rect 27160 27406 27212 27412
rect 26514 27367 26570 27376
rect 26792 26988 26844 26994
rect 26792 26930 26844 26936
rect 26424 26852 26476 26858
rect 26424 26794 26476 26800
rect 26804 26586 26832 26930
rect 27172 26926 27200 27406
rect 27160 26920 27212 26926
rect 27160 26862 27212 26868
rect 27068 26784 27120 26790
rect 27068 26726 27120 26732
rect 25964 26580 26016 26586
rect 25964 26522 26016 26528
rect 26792 26580 26844 26586
rect 26792 26522 26844 26528
rect 25976 26450 26004 26522
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 26240 26376 26292 26382
rect 26240 26318 26292 26324
rect 26252 26042 26280 26318
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26252 25906 26280 25978
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 25516 25498 25544 25842
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 26252 25294 26280 25842
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 24952 24608 25004 24614
rect 24952 24550 25004 24556
rect 24860 24132 24912 24138
rect 24860 24074 24912 24080
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24308 23656 24360 23662
rect 24308 23598 24360 23604
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 24320 23322 24348 23598
rect 24308 23316 24360 23322
rect 24308 23258 24360 23264
rect 24596 23254 24624 23598
rect 24584 23248 24636 23254
rect 24584 23190 24636 23196
rect 24596 22642 24624 23190
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 24308 22432 24360 22438
rect 24308 22374 24360 22380
rect 24320 21554 24348 22374
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24596 21486 24624 22578
rect 24584 21480 24636 21486
rect 24584 21422 24636 21428
rect 24596 21146 24624 21422
rect 24688 21418 24716 22578
rect 24872 21962 24900 24074
rect 24964 23730 24992 24550
rect 24952 23724 25004 23730
rect 24952 23666 25004 23672
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 24964 23118 24992 23666
rect 25700 23526 25728 23666
rect 25688 23520 25740 23526
rect 25688 23462 25740 23468
rect 25792 23186 25820 23666
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 25780 23044 25832 23050
rect 25976 23032 26004 23666
rect 26804 23594 26832 26522
rect 27080 26042 27108 26726
rect 27068 26036 27120 26042
rect 27068 25978 27120 25984
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 27540 23866 27568 25978
rect 27632 25362 27660 28358
rect 27988 27940 28040 27946
rect 27988 27882 28040 27888
rect 28000 25906 28028 27882
rect 28368 27010 28396 31758
rect 28644 31754 28672 32166
rect 29196 31890 29224 32234
rect 29288 31958 29316 32422
rect 29564 32026 29592 32506
rect 29552 32020 29604 32026
rect 29552 31962 29604 31968
rect 29276 31952 29328 31958
rect 29276 31894 29328 31900
rect 29564 31890 29592 31962
rect 29184 31884 29236 31890
rect 29184 31826 29236 31832
rect 29552 31884 29604 31890
rect 29552 31826 29604 31832
rect 29748 31822 29776 32506
rect 30288 32292 30340 32298
rect 30288 32234 30340 32240
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 29000 31816 29052 31822
rect 29000 31758 29052 31764
rect 29736 31816 29788 31822
rect 29736 31758 29788 31764
rect 28644 31726 28764 31754
rect 28448 31204 28500 31210
rect 28448 31146 28500 31152
rect 28460 30734 28488 31146
rect 28448 30728 28500 30734
rect 28448 30670 28500 30676
rect 28736 28966 28764 31726
rect 28816 31748 28868 31754
rect 28816 31690 28868 31696
rect 28828 30734 28856 31690
rect 28908 31680 28960 31686
rect 28908 31622 28960 31628
rect 28920 31278 28948 31622
rect 29012 31328 29040 31758
rect 29748 31346 29776 31758
rect 30116 31754 30144 31826
rect 30104 31748 30156 31754
rect 30104 31690 30156 31696
rect 30116 31346 30144 31690
rect 30300 31346 30328 32234
rect 29092 31340 29144 31346
rect 29012 31300 29092 31328
rect 28908 31272 28960 31278
rect 28908 31214 28960 31220
rect 28920 30938 28948 31214
rect 28908 30932 28960 30938
rect 28908 30874 28960 30880
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 29012 30666 29040 31300
rect 29092 31282 29144 31288
rect 29736 31340 29788 31346
rect 29736 31282 29788 31288
rect 30104 31340 30156 31346
rect 30104 31282 30156 31288
rect 30288 31340 30340 31346
rect 30288 31282 30340 31288
rect 29276 31136 29328 31142
rect 29276 31078 29328 31084
rect 29828 31136 29880 31142
rect 29828 31078 29880 31084
rect 29000 30660 29052 30666
rect 29000 30602 29052 30608
rect 29288 30258 29316 31078
rect 29276 30252 29328 30258
rect 29276 30194 29328 30200
rect 29460 30252 29512 30258
rect 29460 30194 29512 30200
rect 29288 29714 29316 30194
rect 29276 29708 29328 29714
rect 29276 29650 29328 29656
rect 28816 29504 28868 29510
rect 28868 29464 28948 29492
rect 28816 29446 28868 29452
rect 28724 28960 28776 28966
rect 28724 28902 28776 28908
rect 28736 28558 28764 28902
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28552 28218 28580 28494
rect 28540 28212 28592 28218
rect 28540 28154 28592 28160
rect 28724 28008 28776 28014
rect 28724 27950 28776 27956
rect 28736 27674 28764 27950
rect 28724 27668 28776 27674
rect 28724 27610 28776 27616
rect 28632 27396 28684 27402
rect 28632 27338 28684 27344
rect 28276 26994 28396 27010
rect 28644 26994 28672 27338
rect 28264 26988 28396 26994
rect 28316 26982 28396 26988
rect 28264 26930 28316 26936
rect 28368 26450 28396 26982
rect 28632 26988 28684 26994
rect 28632 26930 28684 26936
rect 28540 26920 28592 26926
rect 28540 26862 28592 26868
rect 28448 26852 28500 26858
rect 28448 26794 28500 26800
rect 28356 26444 28408 26450
rect 28356 26386 28408 26392
rect 28172 26240 28224 26246
rect 28172 26182 28224 26188
rect 28184 25906 28212 26182
rect 28368 25906 28396 26386
rect 28460 26042 28488 26794
rect 28448 26036 28500 26042
rect 28448 25978 28500 25984
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 28172 25900 28224 25906
rect 28172 25842 28224 25848
rect 28356 25900 28408 25906
rect 28356 25842 28408 25848
rect 27620 25356 27672 25362
rect 27620 25298 27672 25304
rect 27632 24886 27660 25298
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 27620 24880 27672 24886
rect 27620 24822 27672 24828
rect 27816 24818 27844 25094
rect 27804 24812 27856 24818
rect 27804 24754 27856 24760
rect 27816 24138 27844 24754
rect 28368 24750 28396 25842
rect 28552 25294 28580 26862
rect 28644 26586 28672 26930
rect 28632 26580 28684 26586
rect 28632 26522 28684 26528
rect 28736 25770 28764 27610
rect 28920 27470 28948 29464
rect 29472 29306 29500 30194
rect 29840 29646 29868 31078
rect 30012 30048 30064 30054
rect 30012 29990 30064 29996
rect 30024 29714 30052 29990
rect 30012 29708 30064 29714
rect 30012 29650 30064 29656
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29460 29300 29512 29306
rect 29460 29242 29512 29248
rect 29920 29164 29972 29170
rect 29920 29106 29972 29112
rect 29460 28960 29512 28966
rect 29460 28902 29512 28908
rect 29472 28626 29500 28902
rect 29460 28620 29512 28626
rect 29460 28562 29512 28568
rect 29368 28076 29420 28082
rect 29368 28018 29420 28024
rect 29380 27606 29408 28018
rect 29368 27600 29420 27606
rect 29368 27542 29420 27548
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28920 27334 28948 27406
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 28920 26994 28948 27270
rect 28908 26988 28960 26994
rect 28908 26930 28960 26936
rect 29472 26246 29500 28562
rect 29552 28416 29604 28422
rect 29552 28358 29604 28364
rect 29564 27878 29592 28358
rect 29932 27946 29960 29106
rect 30392 28082 30420 32778
rect 30852 32434 30880 35866
rect 30944 33590 30972 36110
rect 31772 35086 31800 36654
rect 32312 35692 32364 35698
rect 32312 35634 32364 35640
rect 32128 35556 32180 35562
rect 32128 35498 32180 35504
rect 31760 35080 31812 35086
rect 31760 35022 31812 35028
rect 31116 34400 31168 34406
rect 31116 34342 31168 34348
rect 31024 33992 31076 33998
rect 31024 33934 31076 33940
rect 31036 33590 31064 33934
rect 30932 33584 30984 33590
rect 30932 33526 30984 33532
rect 31024 33584 31076 33590
rect 31024 33526 31076 33532
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 30852 30326 30880 32370
rect 31128 32366 31156 34342
rect 31208 33652 31260 33658
rect 31208 33594 31260 33600
rect 31220 33522 31248 33594
rect 31208 33516 31260 33522
rect 31208 33458 31260 33464
rect 31668 33516 31720 33522
rect 31668 33458 31720 33464
rect 31220 32842 31248 33458
rect 31680 33114 31708 33458
rect 31772 33454 31800 35022
rect 32140 34610 32168 35498
rect 32220 35488 32272 35494
rect 32220 35430 32272 35436
rect 32128 34604 32180 34610
rect 32128 34546 32180 34552
rect 32128 34468 32180 34474
rect 32128 34410 32180 34416
rect 32140 34134 32168 34410
rect 32128 34128 32180 34134
rect 32128 34070 32180 34076
rect 32232 33998 32260 35430
rect 32324 34950 32352 35634
rect 32864 35012 32916 35018
rect 32864 34954 32916 34960
rect 32312 34944 32364 34950
rect 32312 34886 32364 34892
rect 32680 34944 32732 34950
rect 32680 34886 32732 34892
rect 32692 34610 32720 34886
rect 32876 34746 32904 34954
rect 32864 34740 32916 34746
rect 32864 34682 32916 34688
rect 32312 34604 32364 34610
rect 32312 34546 32364 34552
rect 32680 34604 32732 34610
rect 32680 34546 32732 34552
rect 32324 34202 32352 34546
rect 32312 34196 32364 34202
rect 32312 34138 32364 34144
rect 32128 33992 32180 33998
rect 32128 33934 32180 33940
rect 32220 33992 32272 33998
rect 32220 33934 32272 33940
rect 31760 33448 31812 33454
rect 31760 33390 31812 33396
rect 31668 33108 31720 33114
rect 31668 33050 31720 33056
rect 31300 32904 31352 32910
rect 31300 32846 31352 32852
rect 31208 32836 31260 32842
rect 31208 32778 31260 32784
rect 31116 32360 31168 32366
rect 31116 32302 31168 32308
rect 31312 31822 31340 32846
rect 31680 32502 31708 33050
rect 31668 32496 31720 32502
rect 31668 32438 31720 32444
rect 31300 31816 31352 31822
rect 31300 31758 31352 31764
rect 31772 31346 31800 33390
rect 32140 32892 32168 33934
rect 32232 33862 32260 33934
rect 32220 33856 32272 33862
rect 32220 33798 32272 33804
rect 32232 33454 32260 33798
rect 32220 33448 32272 33454
rect 32220 33390 32272 33396
rect 32588 33448 32640 33454
rect 32588 33390 32640 33396
rect 32496 33312 32548 33318
rect 32496 33254 32548 33260
rect 32310 33144 32366 33153
rect 32310 33079 32366 33088
rect 32324 33046 32352 33079
rect 32508 33046 32536 33254
rect 32600 33114 32628 33390
rect 32588 33108 32640 33114
rect 32588 33050 32640 33056
rect 32312 33040 32364 33046
rect 32312 32982 32364 32988
rect 32496 33040 32548 33046
rect 32496 32982 32548 32988
rect 32404 32904 32456 32910
rect 32140 32864 32404 32892
rect 32404 32846 32456 32852
rect 32692 32774 32720 34546
rect 32956 34468 33008 34474
rect 32956 34410 33008 34416
rect 32312 32768 32364 32774
rect 32312 32710 32364 32716
rect 32496 32768 32548 32774
rect 32496 32710 32548 32716
rect 32680 32768 32732 32774
rect 32680 32710 32732 32716
rect 32324 31804 32352 32710
rect 32508 32570 32536 32710
rect 32496 32564 32548 32570
rect 32496 32506 32548 32512
rect 32588 32224 32640 32230
rect 32588 32166 32640 32172
rect 32600 31822 32628 32166
rect 32968 31822 32996 34410
rect 33152 33590 33180 36722
rect 34244 36576 34296 36582
rect 34244 36518 34296 36524
rect 34520 36576 34572 36582
rect 34520 36518 34572 36524
rect 35348 36576 35400 36582
rect 35348 36518 35400 36524
rect 34256 36242 34284 36518
rect 34244 36236 34296 36242
rect 34244 36178 34296 36184
rect 33508 35692 33560 35698
rect 33508 35634 33560 35640
rect 33232 35624 33284 35630
rect 33232 35566 33284 35572
rect 33140 33584 33192 33590
rect 33140 33526 33192 33532
rect 33048 33448 33100 33454
rect 33048 33390 33100 33396
rect 33060 31890 33088 33390
rect 33244 33318 33272 35566
rect 33416 35284 33468 35290
rect 33416 35226 33468 35232
rect 33428 34610 33456 35226
rect 33520 34610 33548 35634
rect 34532 34610 34560 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35360 36394 35388 36518
rect 35268 36366 35388 36394
rect 34980 36168 35032 36174
rect 34980 36110 35032 36116
rect 34992 35698 35020 36110
rect 35268 35698 35296 36366
rect 35452 36174 35480 37062
rect 36004 36786 36032 37606
rect 35992 36780 36044 36786
rect 35992 36722 36044 36728
rect 35624 36644 35676 36650
rect 35624 36586 35676 36592
rect 35440 36168 35492 36174
rect 35440 36110 35492 36116
rect 35452 35698 35480 36110
rect 35636 36106 35664 36586
rect 35808 36576 35860 36582
rect 35808 36518 35860 36524
rect 35624 36100 35676 36106
rect 35624 36042 35676 36048
rect 35636 35698 35664 36042
rect 34980 35692 35032 35698
rect 34980 35634 35032 35640
rect 35256 35692 35308 35698
rect 35256 35634 35308 35640
rect 35440 35692 35492 35698
rect 35440 35634 35492 35640
rect 35624 35692 35676 35698
rect 35624 35634 35676 35640
rect 34704 35488 34756 35494
rect 34704 35430 34756 35436
rect 34716 35086 34744 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34704 35080 34756 35086
rect 34704 35022 34756 35028
rect 34888 35080 34940 35086
rect 34888 35022 34940 35028
rect 34716 34762 34744 35022
rect 34624 34734 34744 34762
rect 34900 34746 34928 35022
rect 34980 34944 35032 34950
rect 34980 34886 35032 34892
rect 35440 34944 35492 34950
rect 35440 34886 35492 34892
rect 34888 34740 34940 34746
rect 34624 34678 34652 34734
rect 34888 34682 34940 34688
rect 34612 34672 34664 34678
rect 34612 34614 34664 34620
rect 34992 34610 35020 34886
rect 33416 34604 33468 34610
rect 33416 34546 33468 34552
rect 33508 34604 33560 34610
rect 33508 34546 33560 34552
rect 34428 34604 34480 34610
rect 34428 34546 34480 34552
rect 34520 34604 34572 34610
rect 34520 34546 34572 34552
rect 34704 34604 34756 34610
rect 34704 34546 34756 34552
rect 34980 34604 35032 34610
rect 34980 34546 35032 34552
rect 35348 34604 35400 34610
rect 35348 34546 35400 34552
rect 33324 34400 33376 34406
rect 33324 34342 33376 34348
rect 33336 33522 33364 34342
rect 33428 34134 33456 34546
rect 33416 34128 33468 34134
rect 33416 34070 33468 34076
rect 33416 33992 33468 33998
rect 33416 33934 33468 33940
rect 33324 33516 33376 33522
rect 33324 33458 33376 33464
rect 33232 33312 33284 33318
rect 33232 33254 33284 33260
rect 33138 33144 33194 33153
rect 33138 33079 33140 33088
rect 33192 33079 33194 33088
rect 33140 33050 33192 33056
rect 33244 32910 33272 33254
rect 33232 32904 33284 32910
rect 33232 32846 33284 32852
rect 33140 32836 33192 32842
rect 33140 32778 33192 32784
rect 33152 32570 33180 32778
rect 33140 32564 33192 32570
rect 33140 32506 33192 32512
rect 33336 32502 33364 33458
rect 33428 32910 33456 33934
rect 33520 33522 33548 34546
rect 33968 34536 34020 34542
rect 33968 34478 34020 34484
rect 34440 34490 34468 34546
rect 33980 33998 34008 34478
rect 34440 34462 34560 34490
rect 33968 33992 34020 33998
rect 33968 33934 34020 33940
rect 34532 33930 34560 34462
rect 34716 33998 34744 34546
rect 34796 34400 34848 34406
rect 34796 34342 34848 34348
rect 34704 33992 34756 33998
rect 34704 33934 34756 33940
rect 34428 33924 34480 33930
rect 34428 33866 34480 33872
rect 34520 33924 34572 33930
rect 34520 33866 34572 33872
rect 34440 33522 34468 33866
rect 34808 33522 34836 34342
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 33930 35388 34546
rect 34888 33924 34940 33930
rect 34888 33866 34940 33872
rect 35348 33924 35400 33930
rect 35348 33866 35400 33872
rect 33508 33516 33560 33522
rect 33508 33458 33560 33464
rect 33876 33516 33928 33522
rect 33876 33458 33928 33464
rect 34428 33516 34480 33522
rect 34428 33458 34480 33464
rect 34796 33516 34848 33522
rect 34796 33458 34848 33464
rect 33416 32904 33468 32910
rect 33416 32846 33468 32852
rect 33428 32502 33456 32846
rect 33324 32496 33376 32502
rect 33324 32438 33376 32444
rect 33416 32496 33468 32502
rect 33416 32438 33468 32444
rect 33048 31884 33100 31890
rect 33048 31826 33100 31832
rect 32404 31816 32456 31822
rect 32324 31776 32404 31804
rect 32404 31758 32456 31764
rect 32588 31816 32640 31822
rect 32588 31758 32640 31764
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 33140 31816 33192 31822
rect 33140 31758 33192 31764
rect 32220 31680 32272 31686
rect 32220 31622 32272 31628
rect 31760 31340 31812 31346
rect 31760 31282 31812 31288
rect 32036 31272 32088 31278
rect 32036 31214 32088 31220
rect 30840 30320 30892 30326
rect 30840 30262 30892 30268
rect 30932 29504 30984 29510
rect 30932 29446 30984 29452
rect 31484 29504 31536 29510
rect 32048 29492 32076 31214
rect 32232 30734 32260 31622
rect 33152 30802 33180 31758
rect 33520 31142 33548 33458
rect 33888 32230 33916 33458
rect 34336 33040 34388 33046
rect 34336 32982 34388 32988
rect 34348 32502 34376 32982
rect 34440 32570 34468 33458
rect 34900 33402 34928 33866
rect 35072 33856 35124 33862
rect 35072 33798 35124 33804
rect 35084 33658 35112 33798
rect 35072 33652 35124 33658
rect 35072 33594 35124 33600
rect 34808 33374 34928 33402
rect 34428 32564 34480 32570
rect 34428 32506 34480 32512
rect 34152 32496 34204 32502
rect 34152 32438 34204 32444
rect 34336 32496 34388 32502
rect 34336 32438 34388 32444
rect 33876 32224 33928 32230
rect 33876 32166 33928 32172
rect 33784 31952 33836 31958
rect 33784 31894 33836 31900
rect 33796 31414 33824 31894
rect 34164 31754 34192 32438
rect 34440 31822 34468 32506
rect 34704 31884 34756 31890
rect 34704 31826 34756 31832
rect 34428 31816 34480 31822
rect 34428 31758 34480 31764
rect 34152 31748 34204 31754
rect 34152 31690 34204 31696
rect 33968 31680 34020 31686
rect 33968 31622 34020 31628
rect 33784 31408 33836 31414
rect 33784 31350 33836 31356
rect 33508 31136 33560 31142
rect 33508 31078 33560 31084
rect 33980 30938 34008 31622
rect 33968 30932 34020 30938
rect 33888 30892 33968 30920
rect 33140 30796 33192 30802
rect 33140 30738 33192 30744
rect 32128 30728 32180 30734
rect 32128 30670 32180 30676
rect 32220 30728 32272 30734
rect 32220 30670 32272 30676
rect 32140 29646 32168 30670
rect 33508 30592 33560 30598
rect 33508 30534 33560 30540
rect 33416 30116 33468 30122
rect 33416 30058 33468 30064
rect 32956 29708 33008 29714
rect 32956 29650 33008 29656
rect 32128 29640 32180 29646
rect 32128 29582 32180 29588
rect 32128 29504 32180 29510
rect 32048 29464 32128 29492
rect 31484 29446 31536 29452
rect 32128 29446 32180 29452
rect 30944 29170 30972 29446
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 31496 28082 31524 29446
rect 32140 29238 32168 29446
rect 32128 29232 32180 29238
rect 32128 29174 32180 29180
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31772 28218 31800 29106
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31944 28144 31996 28150
rect 31942 28112 31944 28121
rect 31996 28112 31998 28121
rect 30380 28076 30432 28082
rect 30380 28018 30432 28024
rect 31484 28076 31536 28082
rect 31484 28018 31536 28024
rect 31852 28076 31904 28082
rect 31942 28047 31998 28056
rect 31852 28018 31904 28024
rect 29920 27940 29972 27946
rect 29920 27882 29972 27888
rect 29552 27872 29604 27878
rect 29552 27814 29604 27820
rect 31116 27872 31168 27878
rect 31116 27814 31168 27820
rect 29460 26240 29512 26246
rect 29460 26182 29512 26188
rect 28828 25906 29040 25922
rect 28828 25900 29052 25906
rect 28828 25894 29000 25900
rect 28724 25764 28776 25770
rect 28724 25706 28776 25712
rect 28736 25430 28764 25706
rect 28724 25424 28776 25430
rect 28724 25366 28776 25372
rect 28540 25288 28592 25294
rect 28540 25230 28592 25236
rect 28724 25288 28776 25294
rect 28828 25242 28856 25894
rect 29000 25842 29052 25848
rect 28908 25832 28960 25838
rect 28908 25774 28960 25780
rect 29092 25832 29144 25838
rect 29092 25774 29144 25780
rect 28920 25702 28948 25774
rect 28908 25696 28960 25702
rect 28908 25638 28960 25644
rect 28920 25294 28948 25638
rect 29104 25498 29132 25774
rect 29472 25702 29500 26182
rect 29460 25696 29512 25702
rect 29460 25638 29512 25644
rect 29092 25492 29144 25498
rect 29092 25434 29144 25440
rect 29472 25294 29500 25638
rect 28776 25236 28856 25242
rect 28724 25230 28856 25236
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 29460 25288 29512 25294
rect 29460 25230 29512 25236
rect 28736 25214 28856 25230
rect 28632 25152 28684 25158
rect 28632 25094 28684 25100
rect 28644 24818 28672 25094
rect 28736 24954 28764 25214
rect 29564 25106 29592 27814
rect 30562 27432 30618 27441
rect 31128 27402 31156 27814
rect 30562 27367 30618 27376
rect 31116 27396 31168 27402
rect 29644 26376 29696 26382
rect 29644 26318 29696 26324
rect 29656 25430 29684 26318
rect 29736 26240 29788 26246
rect 29736 26182 29788 26188
rect 29644 25424 29696 25430
rect 29644 25366 29696 25372
rect 29748 25226 29776 26182
rect 30576 25906 30604 27367
rect 31116 27338 31168 27344
rect 31864 27334 31892 28018
rect 31852 27328 31904 27334
rect 31852 27270 31904 27276
rect 30564 25900 30616 25906
rect 30564 25842 30616 25848
rect 31116 25900 31168 25906
rect 31116 25842 31168 25848
rect 29920 25832 29972 25838
rect 29920 25774 29972 25780
rect 29736 25220 29788 25226
rect 29736 25162 29788 25168
rect 29472 25078 29592 25106
rect 28724 24948 28776 24954
rect 28724 24890 28776 24896
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 28816 24200 28868 24206
rect 28816 24142 28868 24148
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 28724 24132 28776 24138
rect 28724 24074 28776 24080
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 27540 23730 27568 23802
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 26792 23588 26844 23594
rect 26792 23530 26844 23536
rect 26424 23520 26476 23526
rect 26424 23462 26476 23468
rect 25832 23004 26004 23032
rect 25780 22986 25832 22992
rect 25792 22234 25820 22986
rect 26436 22234 26464 23462
rect 26804 23050 26832 23530
rect 26988 23322 27016 23666
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 26792 23044 26844 23050
rect 26792 22986 26844 22992
rect 27172 22982 27200 23666
rect 28000 23186 28028 24006
rect 27988 23180 28040 23186
rect 27988 23122 28040 23128
rect 28736 23118 28764 24074
rect 28828 23118 28856 24142
rect 28724 23112 28776 23118
rect 28724 23054 28776 23060
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 27436 22976 27488 22982
rect 27436 22918 27488 22924
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 26424 22228 26476 22234
rect 26424 22170 26476 22176
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 25792 21962 25820 22170
rect 24768 21956 24820 21962
rect 24768 21898 24820 21904
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 25780 21956 25832 21962
rect 25780 21898 25832 21904
rect 24780 21690 24808 21898
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24676 21412 24728 21418
rect 24676 21354 24728 21360
rect 24584 21140 24636 21146
rect 24584 21082 24636 21088
rect 24872 20874 24900 21898
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 26700 21888 26752 21894
rect 26700 21830 26752 21836
rect 26436 21486 26464 21830
rect 26620 21554 26648 21830
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26424 21480 26476 21486
rect 26424 21422 26476 21428
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26252 20942 26280 21286
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24872 19922 24900 20810
rect 26240 20800 26292 20806
rect 26240 20742 26292 20748
rect 26252 20466 26280 20742
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 25884 19786 25912 20198
rect 26344 20058 26372 20402
rect 26436 20330 26464 21422
rect 26712 20942 26740 21830
rect 26988 21486 27016 22170
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 26976 21480 27028 21486
rect 26976 21422 27028 21428
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 26988 20466 27016 21422
rect 27172 21350 27200 21966
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27356 21622 27384 21830
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 27344 20936 27396 20942
rect 27448 20924 27476 22918
rect 27620 22092 27672 22098
rect 27620 22034 27672 22040
rect 28356 22092 28408 22098
rect 28356 22034 28408 22040
rect 27632 21078 27660 22034
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 28000 21146 28028 21286
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 27620 21072 27672 21078
rect 27620 21014 27672 21020
rect 27396 20896 27476 20924
rect 27344 20878 27396 20884
rect 27068 20800 27120 20806
rect 27068 20742 27120 20748
rect 26976 20460 27028 20466
rect 26976 20402 27028 20408
rect 26424 20324 26476 20330
rect 26424 20266 26476 20272
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 27080 19378 27108 20742
rect 27356 20534 27384 20878
rect 28276 20534 28304 21490
rect 27344 20528 27396 20534
rect 27344 20470 27396 20476
rect 28264 20528 28316 20534
rect 28264 20470 28316 20476
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 27160 19780 27212 19786
rect 27160 19722 27212 19728
rect 27172 19514 27200 19722
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 27264 19378 27292 20266
rect 27356 20058 27384 20470
rect 28276 20262 28304 20470
rect 28368 20398 28396 22034
rect 28828 21690 28856 23054
rect 29368 22094 29420 22098
rect 29472 22094 29500 25078
rect 29932 24750 29960 25774
rect 31128 25498 31156 25842
rect 31300 25696 31352 25702
rect 31300 25638 31352 25644
rect 31116 25492 31168 25498
rect 31116 25434 31168 25440
rect 30380 25424 30432 25430
rect 30380 25366 30432 25372
rect 29920 24744 29972 24750
rect 29920 24686 29972 24692
rect 30392 23866 30420 25366
rect 31312 25226 31340 25638
rect 31300 25220 31352 25226
rect 31300 25162 31352 25168
rect 31852 24608 31904 24614
rect 31852 24550 31904 24556
rect 31116 24268 31168 24274
rect 31116 24210 31168 24216
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30380 23860 30432 23866
rect 30380 23802 30432 23808
rect 29552 23520 29604 23526
rect 29552 23462 29604 23468
rect 30012 23520 30064 23526
rect 30012 23462 30064 23468
rect 29564 22642 29592 23462
rect 30024 23186 30052 23462
rect 30012 23180 30064 23186
rect 30012 23122 30064 23128
rect 30288 23044 30340 23050
rect 30288 22986 30340 22992
rect 30300 22710 30328 22986
rect 30392 22982 30420 23802
rect 30852 23730 30880 24006
rect 31128 23730 31156 24210
rect 31864 24206 31892 24550
rect 32140 24342 32168 29174
rect 32404 28212 32456 28218
rect 32404 28154 32456 28160
rect 32312 28144 32364 28150
rect 32232 28104 32312 28132
rect 32232 27334 32260 28104
rect 32312 28086 32364 28092
rect 32416 28082 32444 28154
rect 32404 28076 32456 28082
rect 32404 28018 32456 28024
rect 32220 27328 32272 27334
rect 32220 27270 32272 27276
rect 32232 24818 32260 27270
rect 32312 26376 32364 26382
rect 32312 26318 32364 26324
rect 32324 25294 32352 26318
rect 32416 25838 32444 28018
rect 32968 27470 32996 29650
rect 33428 29646 33456 30058
rect 33520 29646 33548 30534
rect 33888 29696 33916 30892
rect 33968 30874 34020 30880
rect 33704 29668 33916 29696
rect 33416 29640 33468 29646
rect 33416 29582 33468 29588
rect 33508 29640 33560 29646
rect 33508 29582 33560 29588
rect 33140 29504 33192 29510
rect 33140 29446 33192 29452
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 33600 29504 33652 29510
rect 33600 29446 33652 29452
rect 33152 28490 33180 29446
rect 33244 29306 33272 29446
rect 33232 29300 33284 29306
rect 33232 29242 33284 29248
rect 33612 29238 33640 29446
rect 33600 29232 33652 29238
rect 33600 29174 33652 29180
rect 33704 29170 33732 29668
rect 33784 29572 33836 29578
rect 33784 29514 33836 29520
rect 33692 29164 33744 29170
rect 33692 29106 33744 29112
rect 33508 29096 33560 29102
rect 33508 29038 33560 29044
rect 33520 28626 33548 29038
rect 33692 28688 33744 28694
rect 33692 28630 33744 28636
rect 33508 28620 33560 28626
rect 33508 28562 33560 28568
rect 33140 28484 33192 28490
rect 33140 28426 33192 28432
rect 33152 27878 33180 28426
rect 33324 27940 33376 27946
rect 33324 27882 33376 27888
rect 33140 27872 33192 27878
rect 33140 27814 33192 27820
rect 32956 27464 33008 27470
rect 32956 27406 33008 27412
rect 32968 26994 32996 27406
rect 33140 27328 33192 27334
rect 33140 27270 33192 27276
rect 32956 26988 33008 26994
rect 32956 26930 33008 26936
rect 32680 26852 32732 26858
rect 32680 26794 32732 26800
rect 32404 25832 32456 25838
rect 32404 25774 32456 25780
rect 32692 25770 32720 26794
rect 32864 26784 32916 26790
rect 32864 26726 32916 26732
rect 32876 26314 32904 26726
rect 32968 26382 32996 26930
rect 33152 26926 33180 27270
rect 33140 26920 33192 26926
rect 33140 26862 33192 26868
rect 32956 26376 33008 26382
rect 32956 26318 33008 26324
rect 32864 26308 32916 26314
rect 32864 26250 32916 26256
rect 33152 26246 33180 26862
rect 33140 26240 33192 26246
rect 33140 26182 33192 26188
rect 33140 25900 33192 25906
rect 33140 25842 33192 25848
rect 32680 25764 32732 25770
rect 32680 25706 32732 25712
rect 32312 25288 32364 25294
rect 32312 25230 32364 25236
rect 32220 24812 32272 24818
rect 32220 24754 32272 24760
rect 32128 24336 32180 24342
rect 32128 24278 32180 24284
rect 32324 24274 32352 25230
rect 33152 24342 33180 25842
rect 33336 25498 33364 27882
rect 33416 26512 33468 26518
rect 33416 26454 33468 26460
rect 33428 25974 33456 26454
rect 33416 25968 33468 25974
rect 33416 25910 33468 25916
rect 33520 25820 33548 28562
rect 33704 27946 33732 28630
rect 33692 27940 33744 27946
rect 33692 27882 33744 27888
rect 33692 27464 33744 27470
rect 33692 27406 33744 27412
rect 33704 26518 33732 27406
rect 33692 26512 33744 26518
rect 33692 26454 33744 26460
rect 33428 25792 33548 25820
rect 33600 25832 33652 25838
rect 33324 25492 33376 25498
rect 33324 25434 33376 25440
rect 33140 24336 33192 24342
rect 33140 24278 33192 24284
rect 32312 24268 32364 24274
rect 32312 24210 32364 24216
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 31668 24200 31720 24206
rect 31668 24142 31720 24148
rect 31852 24200 31904 24206
rect 31852 24142 31904 24148
rect 31208 23792 31260 23798
rect 31208 23734 31260 23740
rect 30840 23724 30892 23730
rect 30840 23666 30892 23672
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 31116 23724 31168 23730
rect 31116 23666 31168 23672
rect 30748 23656 30800 23662
rect 30748 23598 30800 23604
rect 30760 23338 30788 23598
rect 30576 23310 30788 23338
rect 30472 23248 30524 23254
rect 30472 23190 30524 23196
rect 30380 22976 30432 22982
rect 30380 22918 30432 22924
rect 30288 22704 30340 22710
rect 30288 22646 30340 22652
rect 29552 22636 29604 22642
rect 29552 22578 29604 22584
rect 29828 22636 29880 22642
rect 29828 22578 29880 22584
rect 29368 22092 29500 22094
rect 29420 22066 29500 22092
rect 29368 22034 29420 22040
rect 28816 21684 28868 21690
rect 28816 21626 28868 21632
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 28460 20602 28488 21490
rect 28632 21344 28684 21350
rect 28632 21286 28684 21292
rect 28644 20874 28672 21286
rect 28828 21146 28856 21626
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28632 20868 28684 20874
rect 28632 20810 28684 20816
rect 28448 20596 28500 20602
rect 28448 20538 28500 20544
rect 28828 20466 28856 21082
rect 29564 21010 29592 22578
rect 29840 22234 29868 22578
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30392 21690 30420 22170
rect 30484 22166 30512 23190
rect 30576 23118 30604 23310
rect 30656 23248 30708 23254
rect 30656 23190 30708 23196
rect 30564 23112 30616 23118
rect 30564 23054 30616 23060
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30472 22160 30524 22166
rect 30472 22102 30524 22108
rect 30576 22030 30604 22918
rect 30668 22778 30696 23190
rect 30656 22772 30708 22778
rect 30656 22714 30708 22720
rect 30760 22094 30788 23310
rect 31036 23118 31064 23666
rect 31220 23118 31248 23734
rect 31024 23112 31076 23118
rect 31024 23054 31076 23060
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31036 22930 31064 23054
rect 31036 22902 31156 22930
rect 31024 22772 31076 22778
rect 31024 22714 31076 22720
rect 31036 22098 31064 22714
rect 31128 22234 31156 22902
rect 31496 22778 31524 24142
rect 31484 22772 31536 22778
rect 31484 22714 31536 22720
rect 31680 22642 31708 24142
rect 32324 23730 32352 24210
rect 33152 24206 33180 24278
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 32772 24064 32824 24070
rect 32772 24006 32824 24012
rect 32784 23798 32812 24006
rect 32772 23792 32824 23798
rect 32772 23734 32824 23740
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32324 23322 32352 23666
rect 32312 23316 32364 23322
rect 32312 23258 32364 23264
rect 31668 22636 31720 22642
rect 31668 22578 31720 22584
rect 31208 22432 31260 22438
rect 31208 22374 31260 22380
rect 31116 22228 31168 22234
rect 31116 22170 31168 22176
rect 31128 22098 31156 22170
rect 30668 22066 30788 22094
rect 31024 22092 31076 22098
rect 30564 22024 30616 22030
rect 30564 21966 30616 21972
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 30576 21622 30604 21966
rect 30668 21622 30696 22066
rect 31024 22034 31076 22040
rect 31116 22092 31168 22098
rect 31116 22034 31168 22040
rect 31128 21622 31156 22034
rect 31220 22030 31248 22374
rect 31680 22094 31708 22578
rect 32324 22574 32352 23258
rect 33152 22778 33180 24142
rect 33336 24138 33364 25434
rect 33428 24750 33456 25792
rect 33600 25774 33652 25780
rect 33612 25702 33640 25774
rect 33600 25696 33652 25702
rect 33600 25638 33652 25644
rect 33416 24744 33468 24750
rect 33416 24686 33468 24692
rect 33324 24132 33376 24138
rect 33324 24074 33376 24080
rect 33428 22778 33456 24686
rect 33612 24206 33640 25638
rect 33692 24948 33744 24954
rect 33692 24890 33744 24896
rect 33704 24410 33732 24890
rect 33692 24404 33744 24410
rect 33692 24346 33744 24352
rect 33600 24200 33652 24206
rect 33600 24142 33652 24148
rect 33612 23866 33640 24142
rect 33600 23860 33652 23866
rect 33600 23802 33652 23808
rect 33140 22772 33192 22778
rect 33140 22714 33192 22720
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 32588 22636 32640 22642
rect 32588 22578 32640 22584
rect 32312 22568 32364 22574
rect 32312 22510 32364 22516
rect 32600 22098 32628 22578
rect 31588 22066 31708 22094
rect 31760 22092 31812 22098
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 30564 21616 30616 21622
rect 30564 21558 30616 21564
rect 30656 21616 30708 21622
rect 30656 21558 30708 21564
rect 31116 21616 31168 21622
rect 31116 21558 31168 21564
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 29552 21004 29604 21010
rect 29552 20946 29604 20952
rect 29920 21004 29972 21010
rect 29920 20946 29972 20952
rect 29932 20466 29960 20946
rect 28816 20460 28868 20466
rect 28816 20402 28868 20408
rect 29920 20460 29972 20466
rect 29920 20402 29972 20408
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 30208 20058 30236 20402
rect 30300 20262 30328 21354
rect 30668 21350 30696 21558
rect 31220 21554 31248 21966
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 30668 20602 30696 21286
rect 30656 20596 30708 20602
rect 30656 20538 30708 20544
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 30196 20052 30248 20058
rect 30196 19994 30248 20000
rect 30300 19854 30328 20198
rect 31036 19990 31064 21286
rect 31220 21010 31248 21490
rect 31588 21146 31616 22066
rect 31760 22034 31812 22040
rect 32588 22092 32640 22098
rect 32588 22034 32640 22040
rect 31576 21140 31628 21146
rect 31576 21082 31628 21088
rect 31208 21004 31260 21010
rect 31208 20946 31260 20952
rect 31772 20942 31800 22034
rect 33324 21072 33376 21078
rect 33324 21014 33376 21020
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31772 20754 31800 20878
rect 31772 20726 31892 20754
rect 31760 20392 31812 20398
rect 31760 20334 31812 20340
rect 31024 19984 31076 19990
rect 31024 19926 31076 19932
rect 31772 19922 31800 20334
rect 31760 19916 31812 19922
rect 31760 19858 31812 19864
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 31772 19446 31800 19858
rect 31864 19854 31892 20726
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 33244 19922 33272 20402
rect 33232 19916 33284 19922
rect 33232 19858 33284 19864
rect 31852 19848 31904 19854
rect 31852 19790 31904 19796
rect 32496 19848 32548 19854
rect 32496 19790 32548 19796
rect 32404 19780 32456 19786
rect 32404 19722 32456 19728
rect 32312 19712 32364 19718
rect 32312 19654 32364 19660
rect 31760 19440 31812 19446
rect 31760 19382 31812 19388
rect 32324 19378 32352 19654
rect 32416 19514 32444 19722
rect 32404 19508 32456 19514
rect 32404 19450 32456 19456
rect 32508 19378 32536 19790
rect 33336 19446 33364 21014
rect 33416 20460 33468 20466
rect 33416 20402 33468 20408
rect 33428 19718 33456 20402
rect 33692 20256 33744 20262
rect 33692 20198 33744 20204
rect 33704 19990 33732 20198
rect 33692 19984 33744 19990
rect 33692 19926 33744 19932
rect 33416 19712 33468 19718
rect 33416 19654 33468 19660
rect 33796 19446 33824 29514
rect 33888 28558 33916 29668
rect 34164 29578 34192 31690
rect 34428 31136 34480 31142
rect 34428 31078 34480 31084
rect 34336 29640 34388 29646
rect 34336 29582 34388 29588
rect 34152 29572 34204 29578
rect 34152 29514 34204 29520
rect 33876 28552 33928 28558
rect 33876 28494 33928 28500
rect 34164 28490 34192 29514
rect 34348 29170 34376 29582
rect 34440 29238 34468 31078
rect 34716 30938 34744 31826
rect 34808 31482 34836 33374
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35452 32026 35480 34886
rect 35820 33318 35848 36518
rect 35992 36032 36044 36038
rect 35992 35974 36044 35980
rect 35900 35012 35952 35018
rect 35900 34954 35952 34960
rect 35912 34746 35940 34954
rect 35900 34740 35952 34746
rect 35900 34682 35952 34688
rect 36004 34610 36032 35974
rect 36096 35578 36124 45426
rect 37476 45354 37504 46446
rect 38108 45960 38160 45966
rect 38108 45902 38160 45908
rect 38120 45490 38148 45902
rect 39960 45558 39988 47398
rect 40604 46918 40632 49200
rect 40592 46912 40644 46918
rect 40592 46854 40644 46860
rect 41420 46912 41472 46918
rect 41420 46854 41472 46860
rect 40684 45824 40736 45830
rect 40684 45766 40736 45772
rect 40696 45626 40724 45766
rect 40684 45620 40736 45626
rect 40684 45562 40736 45568
rect 39948 45552 40000 45558
rect 39948 45494 40000 45500
rect 38108 45484 38160 45490
rect 38108 45426 38160 45432
rect 38016 45416 38068 45422
rect 38016 45358 38068 45364
rect 38292 45416 38344 45422
rect 38292 45358 38344 45364
rect 37464 45348 37516 45354
rect 37464 45290 37516 45296
rect 38028 44402 38056 45358
rect 38304 45082 38332 45358
rect 38292 45076 38344 45082
rect 38292 45018 38344 45024
rect 38292 44872 38344 44878
rect 38292 44814 38344 44820
rect 38304 44742 38332 44814
rect 38292 44736 38344 44742
rect 38292 44678 38344 44684
rect 38016 44396 38068 44402
rect 38016 44338 38068 44344
rect 38200 42220 38252 42226
rect 38200 42162 38252 42168
rect 36728 42152 36780 42158
rect 36728 42094 36780 42100
rect 36452 42016 36504 42022
rect 36452 41958 36504 41964
rect 36464 41546 36492 41958
rect 36740 41818 36768 42094
rect 36728 41812 36780 41818
rect 36728 41754 36780 41760
rect 36452 41540 36504 41546
rect 36452 41482 36504 41488
rect 36740 41414 36768 41754
rect 37648 41608 37700 41614
rect 37648 41550 37700 41556
rect 36556 41386 36768 41414
rect 36556 40934 36584 41386
rect 37660 41206 37688 41550
rect 38108 41472 38160 41478
rect 38108 41414 38160 41420
rect 37372 41200 37424 41206
rect 37372 41142 37424 41148
rect 37648 41200 37700 41206
rect 37648 41142 37700 41148
rect 37004 41132 37056 41138
rect 37004 41074 37056 41080
rect 36544 40928 36596 40934
rect 36544 40870 36596 40876
rect 36728 40928 36780 40934
rect 36728 40870 36780 40876
rect 36358 40488 36414 40497
rect 36358 40423 36414 40432
rect 36372 40390 36400 40423
rect 36556 40390 36584 40870
rect 36634 40624 36690 40633
rect 36740 40594 36768 40870
rect 36634 40559 36690 40568
rect 36728 40588 36780 40594
rect 36648 40526 36676 40559
rect 36728 40530 36780 40536
rect 37016 40526 37044 41074
rect 36636 40520 36688 40526
rect 36636 40462 36688 40468
rect 37004 40520 37056 40526
rect 37004 40462 37056 40468
rect 36360 40384 36412 40390
rect 36360 40326 36412 40332
rect 36544 40384 36596 40390
rect 36544 40326 36596 40332
rect 36648 39574 36676 40462
rect 37384 40458 37412 41142
rect 37556 41132 37608 41138
rect 37556 41074 37608 41080
rect 37464 40928 37516 40934
rect 37464 40870 37516 40876
rect 37372 40452 37424 40458
rect 37372 40394 37424 40400
rect 37476 40390 37504 40870
rect 37568 40730 37596 41074
rect 37556 40724 37608 40730
rect 37556 40666 37608 40672
rect 37648 40656 37700 40662
rect 37646 40624 37648 40633
rect 37700 40624 37702 40633
rect 37646 40559 37702 40568
rect 38120 40526 38148 41414
rect 38212 40526 38240 42162
rect 38108 40520 38160 40526
rect 38200 40520 38252 40526
rect 38108 40462 38160 40468
rect 38198 40488 38200 40497
rect 38252 40488 38254 40497
rect 37556 40452 37608 40458
rect 38198 40423 38254 40432
rect 37556 40394 37608 40400
rect 37464 40384 37516 40390
rect 37464 40326 37516 40332
rect 37568 40186 37596 40394
rect 37556 40180 37608 40186
rect 37556 40122 37608 40128
rect 36636 39568 36688 39574
rect 36636 39510 36688 39516
rect 37096 38888 37148 38894
rect 37096 38830 37148 38836
rect 37832 38888 37884 38894
rect 37832 38830 37884 38836
rect 36452 38208 36504 38214
rect 36452 38150 36504 38156
rect 36464 37874 36492 38150
rect 37108 38010 37136 38830
rect 37188 38344 37240 38350
rect 37188 38286 37240 38292
rect 37096 38004 37148 38010
rect 37096 37946 37148 37952
rect 36452 37868 36504 37874
rect 36452 37810 36504 37816
rect 36268 37664 36320 37670
rect 36268 37606 36320 37612
rect 36280 36786 36308 37606
rect 36452 37392 36504 37398
rect 36452 37334 36504 37340
rect 36464 37262 36492 37334
rect 37108 37262 37136 37946
rect 37200 37874 37228 38286
rect 37188 37868 37240 37874
rect 37188 37810 37240 37816
rect 36452 37256 36504 37262
rect 36452 37198 36504 37204
rect 37096 37256 37148 37262
rect 37096 37198 37148 37204
rect 36360 37120 36412 37126
rect 36912 37120 36964 37126
rect 36412 37080 36492 37108
rect 36360 37062 36412 37068
rect 36268 36780 36320 36786
rect 36268 36722 36320 36728
rect 36280 36650 36308 36722
rect 36268 36644 36320 36650
rect 36268 36586 36320 36592
rect 36280 36174 36308 36586
rect 36464 36242 36492 37080
rect 36912 37062 36964 37068
rect 36924 36922 36952 37062
rect 36912 36916 36964 36922
rect 36912 36858 36964 36864
rect 36452 36236 36504 36242
rect 36452 36178 36504 36184
rect 36268 36168 36320 36174
rect 36268 36110 36320 36116
rect 36464 35766 36492 36178
rect 36924 36174 36952 36858
rect 36912 36168 36964 36174
rect 36912 36110 36964 36116
rect 37004 35828 37056 35834
rect 37004 35770 37056 35776
rect 36452 35760 36504 35766
rect 36452 35702 36504 35708
rect 36096 35550 36768 35578
rect 36176 35080 36228 35086
rect 36176 35022 36228 35028
rect 35992 34604 36044 34610
rect 35992 34546 36044 34552
rect 36188 34202 36216 35022
rect 36176 34196 36228 34202
rect 36176 34138 36228 34144
rect 36360 33992 36412 33998
rect 36360 33934 36412 33940
rect 35808 33312 35860 33318
rect 35808 33254 35860 33260
rect 35820 32910 35848 33254
rect 36372 33114 36400 33934
rect 36360 33108 36412 33114
rect 36360 33050 36412 33056
rect 35900 32972 35952 32978
rect 35900 32914 35952 32920
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 35440 32020 35492 32026
rect 35440 31962 35492 31968
rect 34796 31476 34848 31482
rect 34796 31418 34848 31424
rect 34704 30932 34756 30938
rect 34704 30874 34756 30880
rect 34808 30734 34836 31418
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30728 34848 30734
rect 34848 30676 35020 30682
rect 34796 30670 35020 30676
rect 34808 30666 35020 30670
rect 34808 30660 35032 30666
rect 34808 30654 34980 30660
rect 34808 30605 34836 30654
rect 34980 30602 35032 30608
rect 35452 30258 35480 31962
rect 35912 31890 35940 32914
rect 35992 32836 36044 32842
rect 35992 32778 36044 32784
rect 35900 31884 35952 31890
rect 35900 31826 35952 31832
rect 35440 30252 35492 30258
rect 35440 30194 35492 30200
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35900 29776 35952 29782
rect 35900 29718 35952 29724
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 35348 29640 35400 29646
rect 35348 29582 35400 29588
rect 34428 29232 34480 29238
rect 34428 29174 34480 29180
rect 34336 29164 34388 29170
rect 34336 29106 34388 29112
rect 34428 29096 34480 29102
rect 34428 29038 34480 29044
rect 34244 29028 34296 29034
rect 34244 28970 34296 28976
rect 34256 28490 34284 28970
rect 34440 28966 34468 29038
rect 34428 28960 34480 28966
rect 34428 28902 34480 28908
rect 34152 28484 34204 28490
rect 34152 28426 34204 28432
rect 34244 28484 34296 28490
rect 34244 28426 34296 28432
rect 33876 28076 33928 28082
rect 33876 28018 33928 28024
rect 33888 25702 33916 28018
rect 34256 27674 34284 28426
rect 34440 28218 34468 28902
rect 34716 28694 34744 29582
rect 35360 29306 35388 29582
rect 35348 29300 35400 29306
rect 35348 29242 35400 29248
rect 35912 29238 35940 29718
rect 35900 29232 35952 29238
rect 35900 29174 35952 29180
rect 34796 29164 34848 29170
rect 34796 29106 34848 29112
rect 34808 28762 34836 29106
rect 36004 29102 36032 32778
rect 36372 32434 36400 33050
rect 36452 32496 36504 32502
rect 36452 32438 36504 32444
rect 36360 32428 36412 32434
rect 36360 32370 36412 32376
rect 36176 32360 36228 32366
rect 36176 32302 36228 32308
rect 36188 32026 36216 32302
rect 36176 32020 36228 32026
rect 36176 31962 36228 31968
rect 36188 31414 36216 31962
rect 36464 31414 36492 32438
rect 36636 32360 36688 32366
rect 36636 32302 36688 32308
rect 36648 32026 36676 32302
rect 36636 32020 36688 32026
rect 36636 31962 36688 31968
rect 36544 31816 36596 31822
rect 36544 31758 36596 31764
rect 36176 31408 36228 31414
rect 36176 31350 36228 31356
rect 36452 31408 36504 31414
rect 36452 31350 36504 31356
rect 36268 30592 36320 30598
rect 36268 30534 36320 30540
rect 36084 30048 36136 30054
rect 36084 29990 36136 29996
rect 36096 29646 36124 29990
rect 36084 29640 36136 29646
rect 36084 29582 36136 29588
rect 35992 29096 36044 29102
rect 35992 29038 36044 29044
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28756 34848 28762
rect 34796 28698 34848 28704
rect 34704 28688 34756 28694
rect 34704 28630 34756 28636
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 34612 28416 34664 28422
rect 34612 28358 34664 28364
rect 34428 28212 34480 28218
rect 34428 28154 34480 28160
rect 34244 27668 34296 27674
rect 34244 27610 34296 27616
rect 34624 27606 34652 28358
rect 35912 28218 35940 28494
rect 36004 28490 36032 29038
rect 36176 28960 36228 28966
rect 36176 28902 36228 28908
rect 36188 28490 36216 28902
rect 35992 28484 36044 28490
rect 35992 28426 36044 28432
rect 36176 28484 36228 28490
rect 36176 28426 36228 28432
rect 35900 28212 35952 28218
rect 35900 28154 35952 28160
rect 34704 28076 34756 28082
rect 34704 28018 34756 28024
rect 34612 27600 34664 27606
rect 34612 27542 34664 27548
rect 34428 27532 34480 27538
rect 34428 27474 34480 27480
rect 34440 26790 34468 27474
rect 34716 27470 34744 28018
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 35624 27464 35676 27470
rect 35624 27406 35676 27412
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34716 26738 34744 27406
rect 34888 27396 34940 27402
rect 34888 27338 34940 27344
rect 34900 27146 34928 27338
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 34900 27118 35204 27146
rect 35176 26858 35204 27118
rect 35544 27062 35572 27270
rect 35532 27056 35584 27062
rect 35532 26998 35584 27004
rect 35164 26852 35216 26858
rect 35164 26794 35216 26800
rect 34796 26784 34848 26790
rect 34716 26732 34796 26738
rect 34716 26726 34848 26732
rect 34440 26382 34468 26726
rect 34716 26710 34836 26726
rect 34716 26450 34744 26710
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35636 26518 35664 27406
rect 36280 26518 36308 30534
rect 36556 30258 36584 31758
rect 36740 30376 36768 35550
rect 37016 34950 37044 35770
rect 37372 35488 37424 35494
rect 37372 35430 37424 35436
rect 37004 34944 37056 34950
rect 37004 34886 37056 34892
rect 37280 34944 37332 34950
rect 37280 34886 37332 34892
rect 37292 34610 37320 34886
rect 37384 34610 37412 35430
rect 37004 34604 37056 34610
rect 37004 34546 37056 34552
rect 37280 34604 37332 34610
rect 37280 34546 37332 34552
rect 37372 34604 37424 34610
rect 37372 34546 37424 34552
rect 37016 31890 37044 34546
rect 37292 32910 37320 34546
rect 37280 32904 37332 32910
rect 37280 32846 37332 32852
rect 37096 32564 37148 32570
rect 37096 32506 37148 32512
rect 37004 31884 37056 31890
rect 37004 31826 37056 31832
rect 37108 31822 37136 32506
rect 37648 32360 37700 32366
rect 37648 32302 37700 32308
rect 37660 31958 37688 32302
rect 37280 31952 37332 31958
rect 37280 31894 37332 31900
rect 37648 31952 37700 31958
rect 37648 31894 37700 31900
rect 37096 31816 37148 31822
rect 36912 31794 36964 31800
rect 37096 31758 37148 31764
rect 36912 31736 36964 31742
rect 36924 31346 36952 31736
rect 37004 31680 37056 31686
rect 37004 31622 37056 31628
rect 37016 31482 37044 31622
rect 37004 31476 37056 31482
rect 37004 31418 37056 31424
rect 36912 31340 36964 31346
rect 36912 31282 36964 31288
rect 37188 30660 37240 30666
rect 37188 30602 37240 30608
rect 36740 30348 36952 30376
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 36728 30252 36780 30258
rect 36728 30194 36780 30200
rect 36740 29866 36768 30194
rect 36740 29850 36860 29866
rect 36740 29844 36872 29850
rect 36740 29838 36820 29844
rect 36360 29164 36412 29170
rect 36360 29106 36412 29112
rect 36372 28558 36400 29106
rect 36360 28552 36412 28558
rect 36360 28494 36412 28500
rect 36634 28112 36690 28121
rect 36634 28047 36690 28056
rect 36648 28014 36676 28047
rect 36636 28008 36688 28014
rect 36636 27950 36688 27956
rect 36740 27441 36768 29838
rect 36820 29786 36872 29792
rect 36726 27432 36782 27441
rect 36726 27367 36782 27376
rect 36544 26988 36596 26994
rect 36544 26930 36596 26936
rect 35624 26512 35676 26518
rect 35624 26454 35676 26460
rect 36268 26512 36320 26518
rect 36268 26454 36320 26460
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 34428 26376 34480 26382
rect 34428 26318 34480 26324
rect 34440 26042 34468 26318
rect 34428 26036 34480 26042
rect 34428 25978 34480 25984
rect 33876 25696 33928 25702
rect 33876 25638 33928 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35808 25424 35860 25430
rect 35808 25366 35860 25372
rect 35716 24812 35768 24818
rect 35716 24754 35768 24760
rect 33968 24744 34020 24750
rect 33968 24686 34020 24692
rect 35532 24744 35584 24750
rect 35532 24686 35584 24692
rect 33980 24342 34008 24686
rect 34796 24608 34848 24614
rect 34796 24550 34848 24556
rect 33968 24336 34020 24342
rect 33968 24278 34020 24284
rect 33980 24206 34008 24278
rect 34520 24268 34572 24274
rect 34520 24210 34572 24216
rect 33968 24200 34020 24206
rect 33968 24142 34020 24148
rect 34428 23724 34480 23730
rect 34532 23712 34560 24210
rect 34808 24206 34836 24550
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35440 24268 35492 24274
rect 35440 24210 35492 24216
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 34796 24064 34848 24070
rect 34796 24006 34848 24012
rect 35348 24064 35400 24070
rect 35348 24006 35400 24012
rect 34480 23684 34560 23712
rect 34612 23724 34664 23730
rect 34428 23666 34480 23672
rect 34612 23666 34664 23672
rect 34624 23322 34652 23666
rect 34612 23316 34664 23322
rect 34612 23258 34664 23264
rect 34612 21956 34664 21962
rect 34808 21944 34836 24006
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35360 23118 35388 24006
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35452 22098 35480 24210
rect 35544 23526 35572 24686
rect 35728 23730 35756 24754
rect 35820 24206 35848 25366
rect 35900 25288 35952 25294
rect 35900 25230 35952 25236
rect 35992 25288 36044 25294
rect 35992 25230 36044 25236
rect 35912 24682 35940 25230
rect 35900 24676 35952 24682
rect 35900 24618 35952 24624
rect 35808 24200 35860 24206
rect 35808 24142 35860 24148
rect 36004 23866 36032 25230
rect 36280 24138 36308 26454
rect 36452 26240 36504 26246
rect 36452 26182 36504 26188
rect 36464 25906 36492 26182
rect 36452 25900 36504 25906
rect 36452 25842 36504 25848
rect 36464 25226 36492 25842
rect 36556 25702 36584 26930
rect 36544 25696 36596 25702
rect 36544 25638 36596 25644
rect 36556 25498 36584 25638
rect 36544 25492 36596 25498
rect 36544 25434 36596 25440
rect 36452 25220 36504 25226
rect 36452 25162 36504 25168
rect 36268 24132 36320 24138
rect 36268 24074 36320 24080
rect 36176 24064 36228 24070
rect 36176 24006 36228 24012
rect 35992 23860 36044 23866
rect 35992 23802 36044 23808
rect 35716 23724 35768 23730
rect 35716 23666 35768 23672
rect 35532 23520 35584 23526
rect 35532 23462 35584 23468
rect 35544 23118 35572 23462
rect 35728 23322 35756 23666
rect 35716 23316 35768 23322
rect 35716 23258 35768 23264
rect 35532 23112 35584 23118
rect 35532 23054 35584 23060
rect 35900 22976 35952 22982
rect 35900 22918 35952 22924
rect 35912 22710 35940 22918
rect 35900 22704 35952 22710
rect 35900 22646 35952 22652
rect 36004 22642 36032 23802
rect 36188 23798 36216 24006
rect 36176 23792 36228 23798
rect 36176 23734 36228 23740
rect 36464 23118 36492 25162
rect 36636 23520 36688 23526
rect 36636 23462 36688 23468
rect 36452 23112 36504 23118
rect 36452 23054 36504 23060
rect 36648 22642 36676 23462
rect 36924 23322 36952 30348
rect 37004 29232 37056 29238
rect 37004 29174 37056 29180
rect 37016 28558 37044 29174
rect 37004 28552 37056 28558
rect 37004 28494 37056 28500
rect 37004 27328 37056 27334
rect 37004 27270 37056 27276
rect 37016 26314 37044 27270
rect 37004 26308 37056 26314
rect 37004 26250 37056 26256
rect 37200 24614 37228 30602
rect 37292 30258 37320 31894
rect 37844 31754 37872 38830
rect 38200 38820 38252 38826
rect 38200 38762 38252 38768
rect 38212 38350 38240 38762
rect 38200 38344 38252 38350
rect 38200 38286 38252 38292
rect 37924 34060 37976 34066
rect 37924 34002 37976 34008
rect 37936 32570 37964 34002
rect 38108 33380 38160 33386
rect 38108 33322 38160 33328
rect 38016 32904 38068 32910
rect 38016 32846 38068 32852
rect 37924 32564 37976 32570
rect 37924 32506 37976 32512
rect 38028 31890 38056 32846
rect 38016 31884 38068 31890
rect 38016 31826 38068 31832
rect 37844 31726 37964 31754
rect 37280 30252 37332 30258
rect 37280 30194 37332 30200
rect 37372 30252 37424 30258
rect 37372 30194 37424 30200
rect 37556 30252 37608 30258
rect 37556 30194 37608 30200
rect 37384 29730 37412 30194
rect 37384 29702 37504 29730
rect 37568 29714 37596 30194
rect 37648 30116 37700 30122
rect 37648 30058 37700 30064
rect 37372 29640 37424 29646
rect 37372 29582 37424 29588
rect 37280 29504 37332 29510
rect 37280 29446 37332 29452
rect 37292 29170 37320 29446
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37384 28762 37412 29582
rect 37476 29102 37504 29702
rect 37556 29708 37608 29714
rect 37556 29650 37608 29656
rect 37660 29170 37688 30058
rect 37832 30048 37884 30054
rect 37832 29990 37884 29996
rect 37648 29164 37700 29170
rect 37648 29106 37700 29112
rect 37464 29096 37516 29102
rect 37464 29038 37516 29044
rect 37476 28762 37504 29038
rect 37372 28756 37424 28762
rect 37372 28698 37424 28704
rect 37464 28756 37516 28762
rect 37464 28698 37516 28704
rect 37844 28626 37872 29990
rect 37936 29510 37964 31726
rect 38028 29714 38056 31826
rect 38120 30666 38148 33322
rect 38304 31754 38332 44678
rect 40040 43784 40092 43790
rect 40040 43726 40092 43732
rect 40052 43314 40080 43726
rect 40040 43308 40092 43314
rect 40040 43250 40092 43256
rect 41432 43246 41460 46854
rect 41604 46368 41656 46374
rect 41604 46310 41656 46316
rect 41616 46034 41644 46310
rect 42076 46034 42104 49286
rect 42494 49200 42606 50000
rect 43138 49200 43250 50000
rect 44426 49200 44538 50000
rect 45070 49200 45182 50000
rect 46358 49314 46470 50000
rect 45572 49286 46470 49314
rect 45192 47184 45244 47190
rect 45192 47126 45244 47132
rect 41604 46028 41656 46034
rect 41604 45970 41656 45976
rect 42064 46028 42116 46034
rect 42064 45970 42116 45976
rect 41788 45892 41840 45898
rect 41788 45834 41840 45840
rect 41800 45082 41828 45834
rect 45204 45490 45232 47126
rect 45192 45484 45244 45490
rect 45192 45426 45244 45432
rect 41788 45076 41840 45082
rect 41788 45018 41840 45024
rect 41972 44872 42024 44878
rect 41972 44814 42024 44820
rect 40224 43240 40276 43246
rect 40224 43182 40276 43188
rect 41420 43240 41472 43246
rect 41420 43182 41472 43188
rect 40236 42362 40264 43182
rect 40224 42356 40276 42362
rect 40224 42298 40276 42304
rect 41144 42220 41196 42226
rect 41144 42162 41196 42168
rect 41604 42220 41656 42226
rect 41604 42162 41656 42168
rect 40224 42084 40276 42090
rect 40224 42026 40276 42032
rect 40236 41682 40264 42026
rect 40224 41676 40276 41682
rect 40224 41618 40276 41624
rect 39396 41608 39448 41614
rect 39396 41550 39448 41556
rect 40132 41608 40184 41614
rect 40132 41550 40184 41556
rect 39408 41274 39436 41550
rect 40040 41472 40092 41478
rect 40040 41414 40092 41420
rect 40052 41274 40080 41414
rect 39396 41268 39448 41274
rect 39396 41210 39448 41216
rect 40040 41268 40092 41274
rect 40040 41210 40092 41216
rect 40144 40934 40172 41550
rect 40132 40928 40184 40934
rect 40132 40870 40184 40876
rect 40144 40610 40172 40870
rect 40236 40730 40264 41618
rect 40224 40724 40276 40730
rect 40224 40666 40276 40672
rect 40144 40582 40264 40610
rect 40236 40526 40264 40582
rect 40224 40520 40276 40526
rect 40224 40462 40276 40468
rect 38568 39636 38620 39642
rect 38568 39578 38620 39584
rect 38580 35630 38608 39578
rect 39120 39500 39172 39506
rect 39120 39442 39172 39448
rect 39132 38962 39160 39442
rect 39304 39364 39356 39370
rect 39304 39306 39356 39312
rect 39316 38962 39344 39306
rect 39120 38956 39172 38962
rect 39120 38898 39172 38904
rect 39304 38956 39356 38962
rect 39304 38898 39356 38904
rect 38936 38752 38988 38758
rect 38936 38694 38988 38700
rect 40132 38752 40184 38758
rect 40132 38694 40184 38700
rect 38948 37874 38976 38694
rect 40144 37874 40172 38694
rect 40236 38214 40264 40462
rect 40684 40452 40736 40458
rect 40684 40394 40736 40400
rect 40408 39364 40460 39370
rect 40408 39306 40460 39312
rect 40420 39030 40448 39306
rect 40408 39024 40460 39030
rect 40408 38966 40460 38972
rect 40592 38820 40644 38826
rect 40592 38762 40644 38768
rect 40224 38208 40276 38214
rect 40224 38150 40276 38156
rect 40500 38208 40552 38214
rect 40500 38150 40552 38156
rect 38936 37868 38988 37874
rect 38936 37810 38988 37816
rect 40132 37868 40184 37874
rect 40132 37810 40184 37816
rect 40512 37670 40540 38150
rect 40500 37664 40552 37670
rect 40500 37606 40552 37612
rect 39856 36780 39908 36786
rect 39856 36722 39908 36728
rect 38936 35692 38988 35698
rect 38936 35634 38988 35640
rect 38568 35624 38620 35630
rect 38568 35566 38620 35572
rect 38580 34542 38608 35566
rect 38660 35284 38712 35290
rect 38660 35226 38712 35232
rect 38568 34536 38620 34542
rect 38568 34478 38620 34484
rect 38672 33114 38700 35226
rect 38948 35086 38976 35634
rect 39120 35148 39172 35154
rect 39120 35090 39172 35096
rect 38936 35080 38988 35086
rect 38936 35022 38988 35028
rect 38948 34950 38976 35022
rect 38936 34944 38988 34950
rect 38936 34886 38988 34892
rect 39028 34604 39080 34610
rect 39028 34546 39080 34552
rect 38660 33108 38712 33114
rect 38660 33050 38712 33056
rect 38568 32836 38620 32842
rect 38568 32778 38620 32784
rect 38580 32434 38608 32778
rect 38672 32570 38700 33050
rect 39040 32570 39068 34546
rect 39132 34542 39160 35090
rect 39120 34536 39172 34542
rect 39120 34478 39172 34484
rect 39764 33108 39816 33114
rect 39764 33050 39816 33056
rect 38660 32564 38712 32570
rect 38660 32506 38712 32512
rect 39028 32564 39080 32570
rect 39028 32506 39080 32512
rect 39776 32502 39804 33050
rect 39764 32496 39816 32502
rect 39764 32438 39816 32444
rect 38568 32428 38620 32434
rect 38568 32370 38620 32376
rect 38384 32360 38436 32366
rect 38384 32302 38436 32308
rect 38396 31958 38424 32302
rect 38384 31952 38436 31958
rect 38384 31894 38436 31900
rect 38580 31822 38608 32370
rect 38568 31816 38620 31822
rect 38568 31758 38620 31764
rect 38212 31726 38332 31754
rect 38108 30660 38160 30666
rect 38108 30602 38160 30608
rect 38016 29708 38068 29714
rect 38016 29650 38068 29656
rect 37924 29504 37976 29510
rect 37924 29446 37976 29452
rect 38212 28642 38240 31726
rect 38844 31680 38896 31686
rect 38844 31622 38896 31628
rect 38856 31346 38884 31622
rect 38844 31340 38896 31346
rect 38844 31282 38896 31288
rect 39028 31340 39080 31346
rect 39028 31282 39080 31288
rect 38752 31204 38804 31210
rect 38752 31146 38804 31152
rect 38764 30258 38792 31146
rect 38844 31136 38896 31142
rect 38844 31078 38896 31084
rect 38856 30258 38884 31078
rect 39040 30784 39068 31282
rect 39868 30802 39896 36722
rect 40408 36644 40460 36650
rect 40408 36586 40460 36592
rect 40420 36310 40448 36586
rect 40512 36582 40540 37606
rect 40500 36576 40552 36582
rect 40500 36518 40552 36524
rect 40408 36304 40460 36310
rect 40408 36246 40460 36252
rect 39948 35692 40000 35698
rect 39948 35634 40000 35640
rect 39960 34746 39988 35634
rect 40420 35562 40448 36246
rect 40408 35556 40460 35562
rect 40408 35498 40460 35504
rect 40132 35488 40184 35494
rect 40132 35430 40184 35436
rect 40144 35018 40172 35430
rect 40512 35086 40540 36518
rect 40604 35714 40632 38762
rect 40696 35834 40724 40394
rect 41052 39092 41104 39098
rect 41052 39034 41104 39040
rect 40776 38820 40828 38826
rect 40776 38762 40828 38768
rect 40788 38350 40816 38762
rect 41064 38554 41092 39034
rect 40960 38548 41012 38554
rect 40960 38490 41012 38496
rect 41052 38548 41104 38554
rect 41052 38490 41104 38496
rect 40776 38344 40828 38350
rect 40972 38321 41000 38490
rect 40776 38286 40828 38292
rect 40958 38312 41014 38321
rect 40788 38010 40816 38286
rect 40958 38247 41014 38256
rect 40776 38004 40828 38010
rect 40776 37946 40828 37952
rect 40788 37330 40816 37946
rect 40960 37800 41012 37806
rect 40960 37742 41012 37748
rect 40776 37324 40828 37330
rect 40776 37266 40828 37272
rect 40972 37262 41000 37742
rect 40960 37256 41012 37262
rect 40960 37198 41012 37204
rect 40972 36106 41000 37198
rect 40960 36100 41012 36106
rect 40960 36042 41012 36048
rect 40684 35828 40736 35834
rect 40684 35770 40736 35776
rect 40604 35686 40724 35714
rect 40500 35080 40552 35086
rect 40500 35022 40552 35028
rect 40132 35012 40184 35018
rect 40132 34954 40184 34960
rect 40224 34944 40276 34950
rect 40224 34886 40276 34892
rect 39948 34740 40000 34746
rect 39948 34682 40000 34688
rect 40132 33040 40184 33046
rect 40132 32982 40184 32988
rect 40040 32564 40092 32570
rect 40040 32506 40092 32512
rect 39948 32428 40000 32434
rect 39948 32370 40000 32376
rect 39960 31890 39988 32370
rect 39948 31884 40000 31890
rect 39948 31826 40000 31832
rect 40052 31822 40080 32506
rect 40040 31816 40092 31822
rect 40040 31758 40092 31764
rect 38948 30756 39068 30784
rect 39856 30796 39908 30802
rect 38948 30394 38976 30756
rect 39856 30738 39908 30744
rect 40144 30734 40172 32982
rect 40132 30728 40184 30734
rect 40132 30670 40184 30676
rect 39028 30660 39080 30666
rect 39028 30602 39080 30608
rect 38936 30388 38988 30394
rect 38936 30330 38988 30336
rect 38568 30252 38620 30258
rect 38568 30194 38620 30200
rect 38752 30252 38804 30258
rect 38752 30194 38804 30200
rect 38844 30252 38896 30258
rect 38844 30194 38896 30200
rect 38580 29646 38608 30194
rect 38568 29640 38620 29646
rect 38568 29582 38620 29588
rect 38580 28762 38608 29582
rect 38568 28756 38620 28762
rect 38568 28698 38620 28704
rect 37832 28620 37884 28626
rect 37832 28562 37884 28568
rect 38028 28614 38240 28642
rect 37648 28552 37700 28558
rect 37648 28494 37700 28500
rect 37660 27674 37688 28494
rect 37648 27668 37700 27674
rect 37648 27610 37700 27616
rect 37660 27538 37688 27610
rect 37372 27532 37424 27538
rect 37372 27474 37424 27480
rect 37648 27532 37700 27538
rect 37648 27474 37700 27480
rect 37280 27464 37332 27470
rect 37280 27406 37332 27412
rect 37292 26858 37320 27406
rect 37384 27334 37412 27474
rect 37372 27328 37424 27334
rect 37372 27270 37424 27276
rect 37384 26994 37412 27270
rect 37660 27062 37688 27474
rect 37648 27056 37700 27062
rect 37700 27004 37780 27010
rect 37648 26998 37780 27004
rect 37372 26988 37424 26994
rect 37660 26982 37780 26998
rect 37372 26930 37424 26936
rect 37648 26920 37700 26926
rect 37648 26862 37700 26868
rect 37280 26852 37332 26858
rect 37280 26794 37332 26800
rect 37660 26450 37688 26862
rect 37752 26518 37780 26982
rect 37832 26988 37884 26994
rect 37832 26930 37884 26936
rect 37740 26512 37792 26518
rect 37740 26454 37792 26460
rect 37648 26444 37700 26450
rect 37648 26386 37700 26392
rect 37752 26314 37780 26454
rect 37844 26382 37872 26930
rect 38028 26790 38056 28614
rect 38108 28552 38160 28558
rect 38108 28494 38160 28500
rect 38120 27402 38148 28494
rect 38568 27600 38620 27606
rect 38304 27548 38568 27554
rect 38304 27542 38620 27548
rect 38304 27526 38608 27542
rect 38108 27396 38160 27402
rect 38108 27338 38160 27344
rect 38016 26784 38068 26790
rect 38016 26726 38068 26732
rect 38120 26738 38148 27338
rect 38200 26784 38252 26790
rect 38120 26732 38200 26738
rect 38120 26726 38252 26732
rect 38120 26710 38240 26726
rect 37832 26376 37884 26382
rect 37832 26318 37884 26324
rect 38120 26314 38148 26710
rect 38304 26518 38332 27526
rect 38476 27328 38528 27334
rect 38476 27270 38528 27276
rect 38568 27328 38620 27334
rect 38568 27270 38620 27276
rect 38292 26512 38344 26518
rect 38292 26454 38344 26460
rect 38488 26466 38516 27270
rect 38580 26994 38608 27270
rect 38764 26994 38792 30194
rect 38948 29850 38976 30330
rect 38936 29844 38988 29850
rect 38936 29786 38988 29792
rect 38568 26988 38620 26994
rect 38568 26930 38620 26936
rect 38752 26988 38804 26994
rect 38752 26930 38804 26936
rect 38488 26438 38608 26466
rect 38580 26382 38608 26438
rect 38568 26376 38620 26382
rect 38568 26318 38620 26324
rect 37740 26308 37792 26314
rect 37740 26250 37792 26256
rect 38108 26308 38160 26314
rect 38108 26250 38160 26256
rect 38764 24886 38792 26930
rect 39040 25906 39068 30602
rect 40236 29578 40264 34886
rect 40592 33992 40644 33998
rect 40592 33934 40644 33940
rect 40500 32768 40552 32774
rect 40500 32710 40552 32716
rect 40316 32428 40368 32434
rect 40316 32370 40368 32376
rect 40328 31754 40356 32370
rect 40408 31884 40460 31890
rect 40408 31826 40460 31832
rect 40316 31748 40368 31754
rect 40316 31690 40368 31696
rect 40328 30122 40356 31690
rect 40420 31414 40448 31826
rect 40408 31408 40460 31414
rect 40408 31350 40460 31356
rect 40408 30592 40460 30598
rect 40408 30534 40460 30540
rect 40420 30326 40448 30534
rect 40408 30320 40460 30326
rect 40408 30262 40460 30268
rect 40316 30116 40368 30122
rect 40316 30058 40368 30064
rect 40328 29782 40356 30058
rect 40512 29850 40540 32710
rect 40604 30598 40632 33934
rect 40592 30592 40644 30598
rect 40592 30534 40644 30540
rect 40500 29844 40552 29850
rect 40500 29786 40552 29792
rect 40316 29776 40368 29782
rect 40316 29718 40368 29724
rect 40132 29572 40184 29578
rect 40132 29514 40184 29520
rect 40224 29572 40276 29578
rect 40224 29514 40276 29520
rect 40144 28762 40172 29514
rect 40236 28966 40264 29514
rect 40592 29164 40644 29170
rect 40592 29106 40644 29112
rect 40500 29028 40552 29034
rect 40500 28970 40552 28976
rect 40224 28960 40276 28966
rect 40224 28902 40276 28908
rect 40132 28756 40184 28762
rect 40132 28698 40184 28704
rect 40512 28694 40540 28970
rect 40500 28688 40552 28694
rect 40500 28630 40552 28636
rect 40040 28552 40092 28558
rect 40040 28494 40092 28500
rect 39488 27600 39540 27606
rect 39488 27542 39540 27548
rect 39212 27532 39264 27538
rect 39396 27532 39448 27538
rect 39264 27492 39396 27520
rect 39212 27474 39264 27480
rect 39396 27474 39448 27480
rect 39500 27470 39528 27542
rect 39488 27464 39540 27470
rect 39488 27406 39540 27412
rect 39856 26988 39908 26994
rect 39856 26930 39908 26936
rect 39868 26042 39896 26930
rect 39948 26376 40000 26382
rect 39948 26318 40000 26324
rect 39856 26036 39908 26042
rect 39856 25978 39908 25984
rect 39028 25900 39080 25906
rect 39028 25842 39080 25848
rect 38936 25696 38988 25702
rect 38936 25638 38988 25644
rect 38752 24880 38804 24886
rect 38752 24822 38804 24828
rect 37280 24812 37332 24818
rect 37280 24754 37332 24760
rect 37188 24608 37240 24614
rect 37188 24550 37240 24556
rect 37292 24070 37320 24754
rect 38016 24676 38068 24682
rect 38016 24618 38068 24624
rect 38028 24274 38056 24618
rect 38016 24268 38068 24274
rect 38016 24210 38068 24216
rect 38660 24268 38712 24274
rect 38660 24210 38712 24216
rect 38476 24200 38528 24206
rect 38198 24168 38254 24177
rect 38672 24154 38700 24210
rect 38476 24142 38528 24148
rect 38198 24103 38200 24112
rect 38252 24103 38254 24112
rect 38384 24132 38436 24138
rect 38200 24074 38252 24080
rect 38384 24074 38436 24080
rect 37280 24064 37332 24070
rect 37280 24006 37332 24012
rect 37740 24064 37792 24070
rect 37740 24006 37792 24012
rect 36912 23316 36964 23322
rect 36912 23258 36964 23264
rect 37752 23118 37780 24006
rect 38396 23866 38424 24074
rect 38384 23860 38436 23866
rect 38384 23802 38436 23808
rect 38396 23594 38424 23802
rect 38384 23588 38436 23594
rect 38384 23530 38436 23536
rect 37740 23112 37792 23118
rect 37740 23054 37792 23060
rect 37188 22704 37240 22710
rect 37188 22646 37240 22652
rect 35992 22636 36044 22642
rect 35992 22578 36044 22584
rect 36544 22636 36596 22642
rect 36544 22578 36596 22584
rect 36636 22636 36688 22642
rect 36636 22578 36688 22584
rect 36084 22432 36136 22438
rect 36084 22374 36136 22380
rect 35440 22092 35492 22098
rect 35440 22034 35492 22040
rect 34664 21916 34836 21944
rect 34612 21898 34664 21904
rect 34428 21548 34480 21554
rect 34428 21490 34480 21496
rect 33876 21412 33928 21418
rect 33876 21354 33928 21360
rect 33888 20942 33916 21354
rect 33876 20936 33928 20942
rect 33876 20878 33928 20884
rect 34440 20806 34468 21490
rect 34624 21010 34652 21898
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34612 21004 34664 21010
rect 34612 20946 34664 20952
rect 34796 20936 34848 20942
rect 34796 20878 34848 20884
rect 34980 20936 35032 20942
rect 34980 20878 35032 20884
rect 34428 20800 34480 20806
rect 34428 20742 34480 20748
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 33888 20058 33916 20402
rect 33876 20052 33928 20058
rect 33876 19994 33928 20000
rect 34440 19922 34468 20742
rect 34808 20602 34836 20878
rect 34704 20596 34756 20602
rect 34704 20538 34756 20544
rect 34796 20596 34848 20602
rect 34796 20538 34848 20544
rect 34716 20262 34744 20538
rect 34992 20482 35020 20878
rect 35452 20534 35480 22034
rect 35900 21956 35952 21962
rect 35900 21898 35952 21904
rect 35912 21690 35940 21898
rect 35900 21684 35952 21690
rect 35900 21626 35952 21632
rect 36096 21554 36124 22374
rect 36556 21554 36584 22578
rect 37200 21894 37228 22646
rect 37188 21888 37240 21894
rect 37188 21830 37240 21836
rect 36084 21548 36136 21554
rect 36084 21490 36136 21496
rect 36544 21548 36596 21554
rect 36544 21490 36596 21496
rect 37200 21486 37228 21830
rect 38108 21548 38160 21554
rect 38108 21490 38160 21496
rect 37188 21480 37240 21486
rect 37188 21422 37240 21428
rect 35624 20936 35676 20942
rect 35624 20878 35676 20884
rect 34808 20466 35020 20482
rect 35440 20528 35492 20534
rect 35440 20470 35492 20476
rect 34808 20460 35032 20466
rect 34808 20454 34980 20460
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34428 19916 34480 19922
rect 34428 19858 34480 19864
rect 34440 19514 34468 19858
rect 34716 19786 34744 20198
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 34808 19718 34836 20454
rect 34980 20402 35032 20408
rect 34992 20371 35020 20402
rect 35348 20324 35400 20330
rect 35348 20266 35400 20272
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20058 35388 20266
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 35452 19922 35480 20470
rect 35636 20262 35664 20878
rect 37200 20398 37228 21422
rect 37924 21412 37976 21418
rect 37924 21354 37976 21360
rect 37936 20942 37964 21354
rect 38120 21146 38148 21490
rect 38108 21140 38160 21146
rect 38108 21082 38160 21088
rect 38200 21004 38252 21010
rect 38200 20946 38252 20952
rect 37464 20936 37516 20942
rect 37464 20878 37516 20884
rect 37924 20936 37976 20942
rect 37924 20878 37976 20884
rect 37476 20602 37504 20878
rect 37740 20868 37792 20874
rect 37740 20810 37792 20816
rect 37752 20602 37780 20810
rect 37464 20596 37516 20602
rect 37464 20538 37516 20544
rect 37740 20596 37792 20602
rect 37740 20538 37792 20544
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37188 20392 37240 20398
rect 37188 20334 37240 20340
rect 35624 20256 35676 20262
rect 35624 20198 35676 20204
rect 36360 20256 36412 20262
rect 36360 20198 36412 20204
rect 35440 19916 35492 19922
rect 35440 19858 35492 19864
rect 36372 19854 36400 20198
rect 37476 20058 37504 20402
rect 37464 20052 37516 20058
rect 37464 19994 37516 20000
rect 36360 19848 36412 19854
rect 36360 19790 36412 19796
rect 37188 19780 37240 19786
rect 37188 19722 37240 19728
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 34428 19508 34480 19514
rect 34428 19450 34480 19456
rect 37200 19446 37228 19722
rect 37844 19514 37872 20402
rect 38212 20398 38240 20946
rect 38200 20392 38252 20398
rect 38200 20334 38252 20340
rect 38212 19990 38240 20334
rect 38396 20330 38424 23530
rect 38488 23526 38516 24142
rect 38580 24126 38700 24154
rect 38580 23798 38608 24126
rect 38844 24064 38896 24070
rect 38844 24006 38896 24012
rect 38856 23866 38884 24006
rect 38844 23860 38896 23866
rect 38844 23802 38896 23808
rect 38568 23792 38620 23798
rect 38568 23734 38620 23740
rect 38476 23520 38528 23526
rect 38476 23462 38528 23468
rect 38580 23474 38608 23734
rect 38580 23446 38700 23474
rect 38672 22642 38700 23446
rect 38660 22636 38712 22642
rect 38660 22578 38712 22584
rect 38948 22094 38976 25638
rect 39040 23186 39068 25842
rect 39488 24812 39540 24818
rect 39488 24754 39540 24760
rect 39580 24812 39632 24818
rect 39580 24754 39632 24760
rect 39120 24744 39172 24750
rect 39120 24686 39172 24692
rect 39132 24410 39160 24686
rect 39396 24608 39448 24614
rect 39396 24550 39448 24556
rect 39120 24404 39172 24410
rect 39120 24346 39172 24352
rect 39408 24274 39436 24550
rect 39500 24410 39528 24754
rect 39488 24404 39540 24410
rect 39488 24346 39540 24352
rect 39396 24268 39448 24274
rect 39396 24210 39448 24216
rect 39592 23866 39620 24754
rect 39764 24200 39816 24206
rect 39762 24168 39764 24177
rect 39816 24168 39818 24177
rect 39762 24103 39818 24112
rect 39580 23860 39632 23866
rect 39580 23802 39632 23808
rect 39868 23730 39896 25978
rect 39960 25702 39988 26318
rect 39948 25696 40000 25702
rect 39948 25638 40000 25644
rect 40052 24342 40080 28494
rect 40604 28218 40632 29106
rect 40696 28558 40724 35686
rect 40868 35692 40920 35698
rect 40868 35634 40920 35640
rect 40880 34202 40908 35634
rect 40868 34196 40920 34202
rect 40868 34138 40920 34144
rect 40776 33108 40828 33114
rect 40776 33050 40828 33056
rect 40788 29034 40816 33050
rect 40972 32842 41000 36042
rect 41156 34610 41184 42162
rect 41616 41070 41644 42162
rect 41880 42016 41932 42022
rect 41880 41958 41932 41964
rect 41696 41540 41748 41546
rect 41696 41482 41748 41488
rect 41708 41274 41736 41482
rect 41696 41268 41748 41274
rect 41696 41210 41748 41216
rect 41892 41138 41920 41958
rect 41880 41132 41932 41138
rect 41880 41074 41932 41080
rect 41604 41064 41656 41070
rect 41604 41006 41656 41012
rect 41236 40928 41288 40934
rect 41236 40870 41288 40876
rect 41248 40390 41276 40870
rect 41616 40730 41644 41006
rect 41604 40724 41656 40730
rect 41604 40666 41656 40672
rect 41236 40384 41288 40390
rect 41236 40326 41288 40332
rect 41880 39092 41932 39098
rect 41880 39034 41932 39040
rect 41420 39024 41472 39030
rect 41420 38966 41472 38972
rect 41432 38758 41460 38966
rect 41788 38820 41840 38826
rect 41788 38762 41840 38768
rect 41420 38752 41472 38758
rect 41420 38694 41472 38700
rect 41432 37874 41460 38694
rect 41604 38548 41656 38554
rect 41604 38490 41656 38496
rect 41512 38276 41564 38282
rect 41512 38218 41564 38224
rect 41420 37868 41472 37874
rect 41420 37810 41472 37816
rect 41524 37466 41552 38218
rect 41616 38214 41644 38490
rect 41604 38208 41656 38214
rect 41604 38150 41656 38156
rect 41800 38010 41828 38762
rect 41892 38282 41920 39034
rect 41880 38276 41932 38282
rect 41880 38218 41932 38224
rect 41788 38004 41840 38010
rect 41788 37946 41840 37952
rect 41512 37460 41564 37466
rect 41512 37402 41564 37408
rect 41892 37398 41920 38218
rect 41880 37392 41932 37398
rect 41880 37334 41932 37340
rect 41420 37120 41472 37126
rect 41420 37062 41472 37068
rect 41432 36786 41460 37062
rect 41420 36780 41472 36786
rect 41420 36722 41472 36728
rect 41236 36576 41288 36582
rect 41236 36518 41288 36524
rect 41248 36106 41276 36518
rect 41236 36100 41288 36106
rect 41236 36042 41288 36048
rect 41144 34604 41196 34610
rect 41144 34546 41196 34552
rect 40960 32836 41012 32842
rect 40960 32778 41012 32784
rect 40972 32570 41000 32778
rect 40960 32564 41012 32570
rect 40960 32506 41012 32512
rect 41156 31754 41184 34546
rect 41696 34536 41748 34542
rect 41696 34478 41748 34484
rect 41708 34066 41736 34478
rect 41696 34060 41748 34066
rect 41696 34002 41748 34008
rect 41236 33992 41288 33998
rect 41236 33934 41288 33940
rect 41248 33658 41276 33934
rect 41236 33652 41288 33658
rect 41236 33594 41288 33600
rect 41420 33516 41472 33522
rect 41420 33458 41472 33464
rect 41432 33114 41460 33458
rect 41420 33108 41472 33114
rect 41420 33050 41472 33056
rect 41696 33040 41748 33046
rect 41696 32982 41748 32988
rect 41604 32836 41656 32842
rect 41604 32778 41656 32784
rect 41420 31816 41472 31822
rect 41420 31758 41472 31764
rect 40972 31726 41184 31754
rect 40776 29028 40828 29034
rect 40776 28970 40828 28976
rect 40684 28552 40736 28558
rect 40684 28494 40736 28500
rect 40868 28552 40920 28558
rect 40868 28494 40920 28500
rect 40592 28212 40644 28218
rect 40592 28154 40644 28160
rect 40224 28076 40276 28082
rect 40224 28018 40276 28024
rect 40776 28076 40828 28082
rect 40776 28018 40828 28024
rect 40236 26382 40264 28018
rect 40592 27872 40644 27878
rect 40592 27814 40644 27820
rect 40316 27396 40368 27402
rect 40316 27338 40368 27344
rect 40224 26376 40276 26382
rect 40224 26318 40276 26324
rect 40328 25498 40356 27338
rect 40408 26988 40460 26994
rect 40408 26930 40460 26936
rect 40420 26586 40448 26930
rect 40408 26580 40460 26586
rect 40408 26522 40460 26528
rect 40604 26382 40632 27814
rect 40788 27334 40816 28018
rect 40880 27402 40908 28494
rect 40868 27396 40920 27402
rect 40868 27338 40920 27344
rect 40776 27328 40828 27334
rect 40776 27270 40828 27276
rect 40684 26988 40736 26994
rect 40684 26930 40736 26936
rect 40592 26376 40644 26382
rect 40592 26318 40644 26324
rect 40316 25492 40368 25498
rect 40316 25434 40368 25440
rect 40592 24608 40644 24614
rect 40592 24550 40644 24556
rect 40040 24336 40092 24342
rect 40040 24278 40092 24284
rect 39856 23724 39908 23730
rect 39856 23666 39908 23672
rect 40052 23662 40080 24278
rect 40604 23730 40632 24550
rect 40592 23724 40644 23730
rect 40592 23666 40644 23672
rect 40040 23656 40092 23662
rect 40040 23598 40092 23604
rect 39856 23520 39908 23526
rect 39856 23462 39908 23468
rect 39764 23248 39816 23254
rect 39764 23190 39816 23196
rect 39028 23180 39080 23186
rect 39028 23122 39080 23128
rect 39488 22976 39540 22982
rect 39488 22918 39540 22924
rect 39580 22976 39632 22982
rect 39580 22918 39632 22924
rect 39500 22710 39528 22918
rect 39488 22704 39540 22710
rect 39488 22646 39540 22652
rect 39120 22432 39172 22438
rect 39120 22374 39172 22380
rect 39132 22234 39160 22374
rect 39120 22228 39172 22234
rect 39120 22170 39172 22176
rect 38948 22066 39068 22094
rect 38660 21548 38712 21554
rect 38660 21490 38712 21496
rect 38844 21548 38896 21554
rect 38844 21490 38896 21496
rect 38568 21480 38620 21486
rect 38568 21422 38620 21428
rect 38580 21350 38608 21422
rect 38568 21344 38620 21350
rect 38568 21286 38620 21292
rect 38580 20874 38608 21286
rect 38568 20868 38620 20874
rect 38568 20810 38620 20816
rect 38672 20806 38700 21490
rect 38856 21010 38884 21490
rect 38844 21004 38896 21010
rect 38844 20946 38896 20952
rect 39040 20942 39068 22066
rect 39592 22030 39620 22918
rect 39776 22574 39804 23190
rect 39868 23118 39896 23462
rect 39856 23112 39908 23118
rect 39856 23054 39908 23060
rect 39948 23112 40000 23118
rect 39948 23054 40000 23060
rect 40592 23112 40644 23118
rect 40696 23100 40724 26930
rect 40788 26586 40816 27270
rect 40776 26580 40828 26586
rect 40776 26522 40828 26528
rect 40972 25294 41000 31726
rect 41236 31680 41288 31686
rect 41236 31622 41288 31628
rect 41248 31414 41276 31622
rect 41236 31408 41288 31414
rect 41236 31350 41288 31356
rect 41144 31340 41196 31346
rect 41144 31282 41196 31288
rect 41156 30734 41184 31282
rect 41432 30938 41460 31758
rect 41420 30932 41472 30938
rect 41420 30874 41472 30880
rect 41616 30802 41644 32778
rect 41708 32434 41736 32982
rect 41696 32428 41748 32434
rect 41696 32370 41748 32376
rect 41708 31890 41736 32370
rect 41696 31884 41748 31890
rect 41696 31826 41748 31832
rect 41984 31754 42012 44814
rect 45376 44260 45428 44266
rect 45376 44202 45428 44208
rect 45192 44192 45244 44198
rect 45192 44134 45244 44140
rect 45204 42226 45232 44134
rect 45284 42560 45336 42566
rect 45284 42502 45336 42508
rect 42524 42220 42576 42226
rect 42524 42162 42576 42168
rect 45192 42220 45244 42226
rect 45192 42162 45244 42168
rect 42536 41818 42564 42162
rect 43260 42016 43312 42022
rect 43260 41958 43312 41964
rect 42524 41812 42576 41818
rect 42524 41754 42576 41760
rect 42536 41206 42564 41754
rect 43272 41546 43300 41958
rect 45296 41614 45324 42502
rect 45388 42294 45416 44202
rect 45376 42288 45428 42294
rect 45376 42230 45428 42236
rect 43996 41608 44048 41614
rect 43996 41550 44048 41556
rect 45100 41608 45152 41614
rect 45100 41550 45152 41556
rect 45284 41608 45336 41614
rect 45284 41550 45336 41556
rect 43260 41540 43312 41546
rect 43260 41482 43312 41488
rect 43812 41472 43864 41478
rect 43812 41414 43864 41420
rect 42984 41268 43036 41274
rect 42984 41210 43036 41216
rect 42524 41200 42576 41206
rect 42524 41142 42576 41148
rect 42536 40526 42564 41142
rect 42800 40928 42852 40934
rect 42800 40870 42852 40876
rect 42524 40520 42576 40526
rect 42524 40462 42576 40468
rect 42524 40384 42576 40390
rect 42524 40326 42576 40332
rect 42536 39438 42564 40326
rect 42812 39506 42840 40870
rect 42996 40594 43024 41210
rect 43824 41138 43852 41414
rect 44008 41138 44036 41550
rect 43812 41132 43864 41138
rect 43812 41074 43864 41080
rect 43996 41132 44048 41138
rect 43996 41074 44048 41080
rect 44088 41132 44140 41138
rect 44088 41074 44140 41080
rect 42984 40588 43036 40594
rect 42984 40530 43036 40536
rect 43824 40526 43852 41074
rect 43812 40520 43864 40526
rect 43812 40462 43864 40468
rect 42984 40384 43036 40390
rect 42984 40326 43036 40332
rect 42800 39500 42852 39506
rect 42800 39442 42852 39448
rect 42996 39438 43024 40326
rect 44008 39982 44036 41074
rect 44100 40186 44128 41074
rect 44180 40384 44232 40390
rect 44180 40326 44232 40332
rect 44088 40180 44140 40186
rect 44088 40122 44140 40128
rect 44192 40118 44220 40326
rect 44732 40180 44784 40186
rect 44732 40122 44784 40128
rect 44180 40112 44232 40118
rect 44180 40054 44232 40060
rect 43996 39976 44048 39982
rect 43996 39918 44048 39924
rect 42524 39432 42576 39438
rect 42524 39374 42576 39380
rect 42984 39432 43036 39438
rect 42984 39374 43036 39380
rect 42340 39364 42392 39370
rect 42340 39306 42392 39312
rect 42156 38752 42208 38758
rect 42156 38694 42208 38700
rect 42064 38548 42116 38554
rect 42168 38536 42196 38694
rect 42352 38554 42380 39306
rect 42708 39296 42760 39302
rect 42708 39238 42760 39244
rect 42720 38962 42748 39238
rect 44008 38962 44036 39918
rect 42708 38956 42760 38962
rect 42708 38898 42760 38904
rect 43996 38956 44048 38962
rect 43996 38898 44048 38904
rect 42116 38508 42196 38536
rect 42340 38548 42392 38554
rect 42064 38490 42116 38496
rect 42340 38490 42392 38496
rect 44008 38434 44036 38898
rect 42064 38412 42116 38418
rect 42064 38354 42116 38360
rect 43916 38406 44036 38434
rect 42076 38214 42104 38354
rect 43916 38350 43944 38406
rect 42800 38344 42852 38350
rect 42800 38286 42852 38292
rect 43904 38344 43956 38350
rect 43904 38286 43956 38292
rect 42064 38208 42116 38214
rect 42064 38150 42116 38156
rect 42248 37392 42300 37398
rect 42248 37334 42300 37340
rect 42260 36378 42288 37334
rect 42248 36372 42300 36378
rect 42248 36314 42300 36320
rect 42812 36174 42840 38286
rect 43812 38276 43864 38282
rect 43812 38218 43864 38224
rect 44088 38276 44140 38282
rect 44088 38218 44140 38224
rect 43824 38010 43852 38218
rect 43812 38004 43864 38010
rect 43812 37946 43864 37952
rect 44100 37398 44128 38218
rect 44272 37868 44324 37874
rect 44272 37810 44324 37816
rect 44088 37392 44140 37398
rect 44088 37334 44140 37340
rect 44284 37262 44312 37810
rect 43996 37256 44048 37262
rect 44272 37256 44324 37262
rect 44048 37216 44128 37244
rect 43996 37198 44048 37204
rect 43812 37188 43864 37194
rect 43812 37130 43864 37136
rect 42800 36168 42852 36174
rect 42800 36110 42852 36116
rect 42812 34610 42840 36110
rect 42984 36100 43036 36106
rect 42984 36042 43036 36048
rect 42996 35834 43024 36042
rect 42984 35828 43036 35834
rect 42984 35770 43036 35776
rect 42984 35692 43036 35698
rect 42984 35634 43036 35640
rect 42996 35290 43024 35634
rect 43720 35624 43772 35630
rect 43720 35566 43772 35572
rect 43444 35488 43496 35494
rect 43444 35430 43496 35436
rect 42984 35284 43036 35290
rect 42984 35226 43036 35232
rect 42800 34604 42852 34610
rect 42800 34546 42852 34552
rect 42812 33522 42840 34546
rect 42892 33992 42944 33998
rect 42892 33934 42944 33940
rect 42904 33590 42932 33934
rect 43260 33924 43312 33930
rect 43260 33866 43312 33872
rect 43272 33658 43300 33866
rect 43260 33652 43312 33658
rect 43260 33594 43312 33600
rect 43456 33590 43484 35430
rect 43732 35154 43760 35566
rect 43720 35148 43772 35154
rect 43720 35090 43772 35096
rect 43824 34678 43852 37130
rect 43996 36644 44048 36650
rect 43996 36586 44048 36592
rect 44008 35766 44036 36586
rect 44100 36038 44128 37216
rect 44272 37198 44324 37204
rect 44744 36854 44772 40122
rect 45112 39642 45140 41550
rect 45572 41414 45600 49286
rect 46358 49200 46470 49286
rect 47002 49314 47114 50000
rect 47002 49286 48084 49314
rect 47002 49200 47114 49286
rect 46754 49056 46810 49065
rect 46754 48991 46810 49000
rect 46388 47048 46440 47054
rect 46388 46990 46440 46996
rect 46400 46646 46428 46990
rect 46572 46980 46624 46986
rect 46572 46922 46624 46928
rect 46388 46640 46440 46646
rect 46388 46582 46440 46588
rect 46584 46510 46612 46922
rect 46768 46510 46796 48991
rect 46848 47116 46900 47122
rect 46848 47058 46900 47064
rect 46860 47025 46888 47058
rect 47124 47048 47176 47054
rect 46846 47016 46902 47025
rect 47124 46990 47176 46996
rect 46846 46951 46902 46960
rect 46572 46504 46624 46510
rect 46572 46446 46624 46452
rect 46756 46504 46808 46510
rect 46756 46446 46808 46452
rect 45652 46368 45704 46374
rect 45652 46310 45704 46316
rect 46846 46336 46902 46345
rect 45664 45558 45692 46310
rect 46846 46271 46902 46280
rect 45652 45552 45704 45558
rect 45652 45494 45704 45500
rect 46860 45422 46888 46271
rect 47136 45830 47164 46990
rect 47216 46572 47268 46578
rect 47216 46514 47268 46520
rect 47228 46170 47256 46514
rect 47216 46164 47268 46170
rect 47216 46106 47268 46112
rect 47124 45824 47176 45830
rect 47124 45766 47176 45772
rect 46848 45416 46900 45422
rect 46848 45358 46900 45364
rect 46480 44804 46532 44810
rect 46480 44746 46532 44752
rect 46492 44538 46520 44746
rect 46480 44532 46532 44538
rect 46480 44474 46532 44480
rect 46020 43784 46072 43790
rect 46020 43726 46072 43732
rect 46032 43314 46060 43726
rect 46572 43716 46624 43722
rect 46572 43658 46624 43664
rect 46584 43450 46612 43658
rect 46572 43444 46624 43450
rect 46572 43386 46624 43392
rect 46020 43308 46072 43314
rect 46020 43250 46072 43256
rect 46480 43308 46532 43314
rect 46480 43250 46532 43256
rect 45744 42696 45796 42702
rect 45744 42638 45796 42644
rect 45756 42265 45784 42638
rect 45742 42256 45798 42265
rect 45742 42191 45798 42200
rect 46296 42016 46348 42022
rect 46296 41958 46348 41964
rect 46308 41682 46336 41958
rect 46296 41676 46348 41682
rect 46296 41618 46348 41624
rect 46020 41472 46072 41478
rect 46020 41414 46072 41420
rect 46492 41414 46520 43250
rect 46846 42936 46902 42945
rect 46846 42871 46902 42880
rect 46860 42158 46888 42871
rect 46848 42152 46900 42158
rect 46848 42094 46900 42100
rect 46940 41540 46992 41546
rect 46940 41482 46992 41488
rect 45572 41386 45692 41414
rect 45100 39636 45152 39642
rect 45100 39578 45152 39584
rect 45560 38752 45612 38758
rect 45560 38694 45612 38700
rect 45100 38344 45152 38350
rect 45100 38286 45152 38292
rect 45112 38214 45140 38286
rect 45100 38208 45152 38214
rect 45100 38150 45152 38156
rect 44732 36848 44784 36854
rect 44732 36790 44784 36796
rect 44180 36644 44232 36650
rect 44180 36586 44232 36592
rect 44088 36032 44140 36038
rect 44088 35974 44140 35980
rect 44100 35834 44128 35974
rect 44088 35828 44140 35834
rect 44088 35770 44140 35776
rect 43996 35760 44048 35766
rect 43996 35702 44048 35708
rect 44192 35630 44220 36586
rect 44364 35760 44416 35766
rect 44364 35702 44416 35708
rect 44180 35624 44232 35630
rect 44180 35566 44232 35572
rect 44180 35080 44232 35086
rect 44180 35022 44232 35028
rect 43812 34672 43864 34678
rect 43812 34614 43864 34620
rect 43824 34202 43852 34614
rect 43812 34196 43864 34202
rect 43812 34138 43864 34144
rect 43996 33992 44048 33998
rect 43996 33934 44048 33940
rect 42892 33584 42944 33590
rect 42892 33526 42944 33532
rect 43444 33584 43496 33590
rect 43444 33526 43496 33532
rect 42800 33516 42852 33522
rect 42800 33458 42852 33464
rect 42812 33114 42840 33458
rect 42800 33108 42852 33114
rect 42800 33050 42852 33056
rect 42432 32428 42484 32434
rect 42432 32370 42484 32376
rect 42340 31816 42392 31822
rect 42340 31758 42392 31764
rect 41892 31726 42012 31754
rect 41604 30796 41656 30802
rect 41604 30738 41656 30744
rect 41144 30728 41196 30734
rect 41144 30670 41196 30676
rect 41420 30728 41472 30734
rect 41420 30670 41472 30676
rect 41432 30326 41460 30670
rect 41604 30388 41656 30394
rect 41604 30330 41656 30336
rect 41420 30320 41472 30326
rect 41420 30262 41472 30268
rect 41616 30122 41644 30330
rect 41604 30116 41656 30122
rect 41604 30058 41656 30064
rect 41144 29640 41196 29646
rect 41144 29582 41196 29588
rect 41156 29306 41184 29582
rect 41144 29300 41196 29306
rect 41144 29242 41196 29248
rect 41236 28212 41288 28218
rect 41236 28154 41288 28160
rect 41144 28076 41196 28082
rect 41144 28018 41196 28024
rect 41156 27674 41184 28018
rect 41144 27668 41196 27674
rect 41144 27610 41196 27616
rect 41248 26858 41276 28154
rect 41512 27872 41564 27878
rect 41512 27814 41564 27820
rect 41524 27402 41552 27814
rect 41512 27396 41564 27402
rect 41512 27338 41564 27344
rect 41616 26994 41644 30058
rect 41604 26988 41656 26994
rect 41604 26930 41656 26936
rect 41236 26852 41288 26858
rect 41236 26794 41288 26800
rect 41248 26450 41276 26794
rect 41236 26444 41288 26450
rect 41236 26386 41288 26392
rect 41604 26308 41656 26314
rect 41604 26250 41656 26256
rect 41616 25906 41644 26250
rect 41892 25974 41920 31726
rect 41972 31136 42024 31142
rect 41972 31078 42024 31084
rect 41984 30802 42012 31078
rect 42352 30938 42380 31758
rect 42340 30932 42392 30938
rect 42340 30874 42392 30880
rect 41972 30796 42024 30802
rect 41972 30738 42024 30744
rect 42444 28014 42472 32370
rect 42800 32020 42852 32026
rect 42800 31962 42852 31968
rect 42524 31952 42576 31958
rect 42524 31894 42576 31900
rect 42536 30258 42564 31894
rect 42812 30802 42840 31962
rect 42904 31754 42932 33526
rect 44008 32910 44036 33934
rect 44192 33114 44220 35022
rect 44180 33108 44232 33114
rect 44180 33050 44232 33056
rect 43996 32904 44048 32910
rect 43996 32846 44048 32852
rect 43536 32428 43588 32434
rect 43536 32370 43588 32376
rect 43352 32360 43404 32366
rect 43352 32302 43404 32308
rect 42904 31726 43024 31754
rect 42892 31476 42944 31482
rect 42892 31418 42944 31424
rect 42904 31346 42932 31418
rect 42892 31340 42944 31346
rect 42892 31282 42944 31288
rect 42800 30796 42852 30802
rect 42800 30738 42852 30744
rect 42524 30252 42576 30258
rect 42524 30194 42576 30200
rect 42996 28490 43024 31726
rect 43168 31680 43220 31686
rect 43168 31622 43220 31628
rect 43076 31272 43128 31278
rect 43076 31214 43128 31220
rect 43088 30734 43116 31214
rect 43180 31142 43208 31622
rect 43364 31482 43392 32302
rect 43548 32026 43576 32370
rect 44180 32224 44232 32230
rect 44180 32166 44232 32172
rect 43536 32020 43588 32026
rect 43536 31962 43588 31968
rect 43444 31816 43496 31822
rect 43444 31758 43496 31764
rect 43352 31476 43404 31482
rect 43352 31418 43404 31424
rect 43168 31136 43220 31142
rect 43168 31078 43220 31084
rect 43076 30728 43128 30734
rect 43076 30670 43128 30676
rect 43456 29850 43484 31758
rect 43628 31748 43680 31754
rect 43628 31690 43680 31696
rect 43640 31414 43668 31690
rect 43904 31680 43956 31686
rect 43904 31622 43956 31628
rect 43996 31680 44048 31686
rect 43996 31622 44048 31628
rect 43628 31408 43680 31414
rect 43628 31350 43680 31356
rect 43916 31346 43944 31622
rect 44008 31482 44036 31622
rect 43996 31476 44048 31482
rect 43996 31418 44048 31424
rect 44192 31414 44220 32166
rect 44272 31680 44324 31686
rect 44272 31622 44324 31628
rect 44180 31408 44232 31414
rect 44180 31350 44232 31356
rect 43904 31340 43956 31346
rect 43904 31282 43956 31288
rect 43812 31272 43864 31278
rect 43812 31214 43864 31220
rect 43824 30326 43852 31214
rect 43812 30320 43864 30326
rect 43812 30262 43864 30268
rect 43824 30190 43852 30262
rect 43812 30184 43864 30190
rect 43812 30126 43864 30132
rect 43444 29844 43496 29850
rect 43444 29786 43496 29792
rect 43456 29730 43484 29786
rect 43364 29702 43484 29730
rect 43260 29572 43312 29578
rect 43260 29514 43312 29520
rect 43272 29050 43300 29514
rect 43364 29170 43392 29702
rect 43444 29640 43496 29646
rect 43444 29582 43496 29588
rect 43456 29306 43484 29582
rect 43444 29300 43496 29306
rect 43444 29242 43496 29248
rect 43352 29164 43404 29170
rect 43352 29106 43404 29112
rect 43824 29102 43852 30126
rect 43916 30054 43944 31282
rect 44180 30864 44232 30870
rect 44180 30806 44232 30812
rect 43904 30048 43956 30054
rect 43904 29990 43956 29996
rect 44192 29238 44220 30806
rect 44284 30802 44312 31622
rect 44376 30802 44404 35702
rect 44640 35692 44692 35698
rect 44640 35634 44692 35640
rect 44652 33674 44680 35634
rect 44744 35494 44772 36790
rect 45112 36564 45140 38150
rect 45572 37874 45600 38694
rect 45560 37868 45612 37874
rect 45560 37810 45612 37816
rect 45192 36576 45244 36582
rect 45112 36536 45192 36564
rect 45192 36518 45244 36524
rect 45204 35630 45232 36518
rect 45572 36242 45600 37810
rect 45560 36236 45612 36242
rect 45560 36178 45612 36184
rect 45192 35624 45244 35630
rect 45192 35566 45244 35572
rect 44732 35488 44784 35494
rect 44732 35430 44784 35436
rect 44744 35086 44772 35430
rect 44732 35080 44784 35086
rect 44732 35022 44784 35028
rect 45192 34944 45244 34950
rect 45192 34886 45244 34892
rect 45008 34604 45060 34610
rect 45008 34546 45060 34552
rect 45020 34202 45048 34546
rect 45008 34196 45060 34202
rect 45008 34138 45060 34144
rect 45204 33998 45232 34886
rect 45192 33992 45244 33998
rect 45192 33934 45244 33940
rect 44560 33646 44680 33674
rect 44456 32428 44508 32434
rect 44456 32370 44508 32376
rect 44468 30938 44496 32370
rect 44456 30932 44508 30938
rect 44456 30874 44508 30880
rect 44272 30796 44324 30802
rect 44272 30738 44324 30744
rect 44364 30796 44416 30802
rect 44364 30738 44416 30744
rect 44456 30728 44508 30734
rect 44456 30670 44508 30676
rect 44468 29510 44496 30670
rect 44272 29504 44324 29510
rect 44272 29446 44324 29452
rect 44456 29504 44508 29510
rect 44456 29446 44508 29452
rect 44180 29232 44232 29238
rect 44180 29174 44232 29180
rect 43812 29096 43864 29102
rect 43272 29022 43392 29050
rect 43812 29038 43864 29044
rect 43364 28558 43392 29022
rect 43352 28552 43404 28558
rect 43352 28494 43404 28500
rect 42984 28484 43036 28490
rect 42984 28426 43036 28432
rect 42432 28008 42484 28014
rect 42432 27950 42484 27956
rect 42616 28008 42668 28014
rect 42616 27950 42668 27956
rect 41880 25968 41932 25974
rect 41880 25910 41932 25916
rect 41604 25900 41656 25906
rect 41604 25842 41656 25848
rect 41604 25356 41656 25362
rect 41604 25298 41656 25304
rect 40960 25288 41012 25294
rect 40960 25230 41012 25236
rect 40972 24954 41000 25230
rect 41420 25152 41472 25158
rect 41420 25094 41472 25100
rect 40960 24948 41012 24954
rect 40960 24890 41012 24896
rect 41432 24274 41460 25094
rect 41420 24268 41472 24274
rect 41420 24210 41472 24216
rect 41236 24200 41288 24206
rect 41236 24142 41288 24148
rect 41248 23322 41276 24142
rect 41144 23316 41196 23322
rect 41144 23258 41196 23264
rect 41236 23316 41288 23322
rect 41236 23258 41288 23264
rect 40644 23072 40724 23100
rect 40592 23054 40644 23060
rect 39960 22710 39988 23054
rect 40040 23044 40092 23050
rect 40040 22986 40092 22992
rect 40052 22778 40080 22986
rect 40132 22976 40184 22982
rect 40132 22918 40184 22924
rect 40040 22772 40092 22778
rect 40040 22714 40092 22720
rect 39948 22704 40000 22710
rect 39948 22646 40000 22652
rect 40144 22642 40172 22918
rect 40132 22636 40184 22642
rect 40132 22578 40184 22584
rect 40316 22636 40368 22642
rect 40316 22578 40368 22584
rect 40408 22636 40460 22642
rect 40408 22578 40460 22584
rect 39764 22568 39816 22574
rect 39684 22528 39764 22556
rect 39580 22024 39632 22030
rect 39580 21966 39632 21972
rect 39488 21888 39540 21894
rect 39488 21830 39540 21836
rect 39500 21554 39528 21830
rect 39488 21548 39540 21554
rect 39488 21490 39540 21496
rect 39120 21072 39172 21078
rect 39120 21014 39172 21020
rect 39028 20936 39080 20942
rect 39028 20878 39080 20884
rect 38660 20800 38712 20806
rect 38660 20742 38712 20748
rect 39132 20466 39160 21014
rect 39592 21010 39620 21966
rect 39580 21004 39632 21010
rect 39580 20946 39632 20952
rect 39304 20936 39356 20942
rect 39304 20878 39356 20884
rect 39316 20602 39344 20878
rect 39488 20800 39540 20806
rect 39488 20742 39540 20748
rect 39304 20596 39356 20602
rect 39304 20538 39356 20544
rect 39120 20460 39172 20466
rect 39120 20402 39172 20408
rect 38384 20324 38436 20330
rect 38384 20266 38436 20272
rect 38200 19984 38252 19990
rect 38200 19926 38252 19932
rect 39316 19922 39344 20538
rect 39500 20466 39528 20742
rect 39488 20460 39540 20466
rect 39488 20402 39540 20408
rect 39304 19916 39356 19922
rect 39304 19858 39356 19864
rect 39684 19854 39712 22528
rect 39764 22510 39816 22516
rect 40328 22234 40356 22578
rect 40420 22438 40448 22578
rect 40592 22568 40644 22574
rect 40592 22510 40644 22516
rect 40408 22432 40460 22438
rect 40408 22374 40460 22380
rect 39856 22228 39908 22234
rect 39856 22170 39908 22176
rect 40316 22228 40368 22234
rect 40316 22170 40368 22176
rect 39868 21962 39896 22170
rect 40420 22030 40448 22374
rect 39948 22024 40000 22030
rect 39948 21966 40000 21972
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 40408 22024 40460 22030
rect 40408 21966 40460 21972
rect 39856 21956 39908 21962
rect 39856 21898 39908 21904
rect 39868 21554 39896 21898
rect 39960 21690 39988 21966
rect 39948 21684 40000 21690
rect 39948 21626 40000 21632
rect 40052 21554 40080 21966
rect 40604 21962 40632 22510
rect 40696 22030 40724 23072
rect 40776 23112 40828 23118
rect 40776 23054 40828 23060
rect 40788 22778 40816 23054
rect 41156 22778 41184 23258
rect 40776 22772 40828 22778
rect 40776 22714 40828 22720
rect 41144 22772 41196 22778
rect 41144 22714 41196 22720
rect 41512 22500 41564 22506
rect 41512 22442 41564 22448
rect 41420 22092 41472 22098
rect 41420 22034 41472 22040
rect 40684 22024 40736 22030
rect 40684 21966 40736 21972
rect 40592 21956 40644 21962
rect 40592 21898 40644 21904
rect 39856 21548 39908 21554
rect 39856 21490 39908 21496
rect 40040 21548 40092 21554
rect 40040 21490 40092 21496
rect 39764 21480 39816 21486
rect 39764 21422 39816 21428
rect 39776 21146 39804 21422
rect 39764 21140 39816 21146
rect 39764 21082 39816 21088
rect 39120 19848 39172 19854
rect 39120 19790 39172 19796
rect 39672 19848 39724 19854
rect 39672 19790 39724 19796
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 37832 19508 37884 19514
rect 37832 19450 37884 19456
rect 33324 19440 33376 19446
rect 33324 19382 33376 19388
rect 33784 19440 33836 19446
rect 33784 19382 33836 19388
rect 37188 19440 37240 19446
rect 37188 19382 37240 19388
rect 27068 19372 27120 19378
rect 27068 19314 27120 19320
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 37844 17678 37872 19450
rect 38752 19372 38804 19378
rect 38752 19314 38804 19320
rect 38764 18902 38792 19314
rect 38856 18970 38884 19654
rect 39132 19378 39160 19790
rect 39120 19372 39172 19378
rect 39120 19314 39172 19320
rect 38844 18964 38896 18970
rect 38844 18906 38896 18912
rect 40052 18902 40080 21490
rect 41432 20874 41460 22034
rect 41420 20868 41472 20874
rect 41420 20810 41472 20816
rect 41524 20058 41552 22442
rect 40500 20052 40552 20058
rect 40500 19994 40552 20000
rect 41512 20052 41564 20058
rect 41512 19994 41564 20000
rect 40224 19848 40276 19854
rect 40224 19790 40276 19796
rect 40236 19446 40264 19790
rect 40316 19780 40368 19786
rect 40316 19722 40368 19728
rect 40224 19440 40276 19446
rect 40224 19382 40276 19388
rect 40328 19378 40356 19722
rect 40316 19372 40368 19378
rect 40316 19314 40368 19320
rect 40408 19372 40460 19378
rect 40512 19360 40540 19994
rect 40868 19712 40920 19718
rect 40868 19654 40920 19660
rect 40776 19440 40828 19446
rect 40776 19382 40828 19388
rect 40460 19332 40540 19360
rect 40408 19314 40460 19320
rect 38752 18896 38804 18902
rect 38752 18838 38804 18844
rect 40040 18896 40092 18902
rect 40040 18838 40092 18844
rect 40408 18760 40460 18766
rect 40408 18702 40460 18708
rect 39212 18692 39264 18698
rect 39212 18634 39264 18640
rect 39224 17814 39252 18634
rect 39212 17808 39264 17814
rect 39212 17750 39264 17756
rect 37832 17672 37884 17678
rect 37832 17614 37884 17620
rect 39856 17672 39908 17678
rect 39856 17614 39908 17620
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 39868 16794 39896 17614
rect 40420 17338 40448 18702
rect 40512 17746 40540 19332
rect 40788 18970 40816 19382
rect 40880 19378 40908 19654
rect 40868 19372 40920 19378
rect 40868 19314 40920 19320
rect 40776 18964 40828 18970
rect 40776 18906 40828 18912
rect 41616 18834 41644 25298
rect 42432 23792 42484 23798
rect 42432 23734 42484 23740
rect 42444 22642 42472 23734
rect 42064 22636 42116 22642
rect 42064 22578 42116 22584
rect 42432 22636 42484 22642
rect 42432 22578 42484 22584
rect 42524 22636 42576 22642
rect 42524 22578 42576 22584
rect 41788 22024 41840 22030
rect 41788 21966 41840 21972
rect 41972 22002 42024 22008
rect 41800 21078 41828 21966
rect 41972 21944 42024 21950
rect 41984 21690 42012 21944
rect 41972 21684 42024 21690
rect 41972 21626 42024 21632
rect 41880 21548 41932 21554
rect 41880 21490 41932 21496
rect 41788 21072 41840 21078
rect 41788 21014 41840 21020
rect 41892 20602 41920 21490
rect 41696 20596 41748 20602
rect 41696 20538 41748 20544
rect 41880 20596 41932 20602
rect 41880 20538 41932 20544
rect 41708 19446 41736 20538
rect 41880 20256 41932 20262
rect 41880 20198 41932 20204
rect 41696 19440 41748 19446
rect 41696 19382 41748 19388
rect 41892 19242 41920 20198
rect 42076 19922 42104 22578
rect 42536 22234 42564 22578
rect 42524 22228 42576 22234
rect 42524 22170 42576 22176
rect 42628 22094 42656 27950
rect 42892 27396 42944 27402
rect 42892 27338 42944 27344
rect 42904 26994 42932 27338
rect 43364 27130 43392 28494
rect 43824 27878 43852 29038
rect 44088 28756 44140 28762
rect 44088 28698 44140 28704
rect 43812 27872 43864 27878
rect 43812 27814 43864 27820
rect 43824 27470 43852 27814
rect 43812 27464 43864 27470
rect 43812 27406 43864 27412
rect 43444 27328 43496 27334
rect 43444 27270 43496 27276
rect 43352 27124 43404 27130
rect 43352 27066 43404 27072
rect 42892 26988 42944 26994
rect 42892 26930 42944 26936
rect 43456 25226 43484 27270
rect 43824 26926 43852 27406
rect 44100 27062 44128 28698
rect 44284 28150 44312 29446
rect 44560 28762 44588 33646
rect 44824 33516 44876 33522
rect 44824 33458 44876 33464
rect 44732 33380 44784 33386
rect 44732 33322 44784 33328
rect 44640 33312 44692 33318
rect 44640 33254 44692 33260
rect 44652 32910 44680 33254
rect 44640 32904 44692 32910
rect 44640 32846 44692 32852
rect 44548 28756 44600 28762
rect 44548 28698 44600 28704
rect 44744 28626 44772 33322
rect 44836 32570 44864 33458
rect 44824 32564 44876 32570
rect 44824 32506 44876 32512
rect 45664 31754 45692 41386
rect 46032 41138 46060 41414
rect 46492 41386 46704 41414
rect 46676 41138 46704 41386
rect 46952 41274 46980 41482
rect 46940 41268 46992 41274
rect 46940 41210 46992 41216
rect 46020 41132 46072 41138
rect 46020 41074 46072 41080
rect 46664 41132 46716 41138
rect 46664 41074 46716 41080
rect 45836 40928 45888 40934
rect 45836 40870 45888 40876
rect 46296 40928 46348 40934
rect 46296 40870 46348 40876
rect 45848 40050 45876 40870
rect 46308 40594 46336 40870
rect 46296 40588 46348 40594
rect 46296 40530 46348 40536
rect 46478 40216 46534 40225
rect 46478 40151 46534 40160
rect 45836 40044 45888 40050
rect 45836 39986 45888 39992
rect 45928 38412 45980 38418
rect 45928 38354 45980 38360
rect 45836 36576 45888 36582
rect 45836 36518 45888 36524
rect 45848 36378 45876 36518
rect 45836 36372 45888 36378
rect 45836 36314 45888 36320
rect 45940 36174 45968 38354
rect 46296 38208 46348 38214
rect 46296 38150 46348 38156
rect 46308 37874 46336 38150
rect 46296 37868 46348 37874
rect 46296 37810 46348 37816
rect 46296 37256 46348 37262
rect 46296 37198 46348 37204
rect 46308 36854 46336 37198
rect 46204 36848 46256 36854
rect 46204 36790 46256 36796
rect 46296 36848 46348 36854
rect 46296 36790 46348 36796
rect 46216 36378 46244 36790
rect 46204 36372 46256 36378
rect 46204 36314 46256 36320
rect 45928 36168 45980 36174
rect 45928 36110 45980 36116
rect 45744 35692 45796 35698
rect 45744 35634 45796 35640
rect 45756 35154 45784 35634
rect 45940 35578 45968 36110
rect 46388 36032 46440 36038
rect 46388 35974 46440 35980
rect 46400 35698 46428 35974
rect 46388 35692 46440 35698
rect 46388 35634 46440 35640
rect 45940 35550 46060 35578
rect 46032 35494 46060 35550
rect 46020 35488 46072 35494
rect 46020 35430 46072 35436
rect 45744 35148 45796 35154
rect 45744 35090 45796 35096
rect 45756 34746 45784 35090
rect 45744 34740 45796 34746
rect 45744 34682 45796 34688
rect 46400 34610 46428 35634
rect 46388 34604 46440 34610
rect 46388 34546 46440 34552
rect 46492 34066 46520 40151
rect 46572 38752 46624 38758
rect 46572 38694 46624 38700
rect 46584 38418 46612 38694
rect 46572 38412 46624 38418
rect 46572 38354 46624 38360
rect 46676 36582 46704 41074
rect 46940 40452 46992 40458
rect 46940 40394 46992 40400
rect 46952 40050 46980 40394
rect 46940 40044 46992 40050
rect 46940 39986 46992 39992
rect 46756 38956 46808 38962
rect 46756 38898 46808 38904
rect 46768 38554 46796 38898
rect 46756 38548 46808 38554
rect 46756 38490 46808 38496
rect 46940 37664 46992 37670
rect 46940 37606 46992 37612
rect 46664 36576 46716 36582
rect 46664 36518 46716 36524
rect 46848 36576 46900 36582
rect 46848 36518 46900 36524
rect 46572 36100 46624 36106
rect 46572 36042 46624 36048
rect 46584 35630 46612 36042
rect 46572 35624 46624 35630
rect 46572 35566 46624 35572
rect 46584 35290 46612 35566
rect 46572 35284 46624 35290
rect 46572 35226 46624 35232
rect 46480 34060 46532 34066
rect 46480 34002 46532 34008
rect 46112 32768 46164 32774
rect 46112 32710 46164 32716
rect 45664 31726 45968 31754
rect 45744 31340 45796 31346
rect 45744 31282 45796 31288
rect 44824 31204 44876 31210
rect 44824 31146 44876 31152
rect 44836 30598 44864 31146
rect 45100 31136 45152 31142
rect 45100 31078 45152 31084
rect 45112 30666 45140 31078
rect 45652 30728 45704 30734
rect 45652 30670 45704 30676
rect 45100 30660 45152 30666
rect 45100 30602 45152 30608
rect 44824 30592 44876 30598
rect 44824 30534 44876 30540
rect 45664 30190 45692 30670
rect 45756 30666 45784 31282
rect 45744 30660 45796 30666
rect 45744 30602 45796 30608
rect 45652 30184 45704 30190
rect 45652 30126 45704 30132
rect 45008 29300 45060 29306
rect 45008 29242 45060 29248
rect 44732 28620 44784 28626
rect 44732 28562 44784 28568
rect 44272 28144 44324 28150
rect 44272 28086 44324 28092
rect 44088 27056 44140 27062
rect 44088 26998 44140 27004
rect 43812 26920 43864 26926
rect 43812 26862 43864 26868
rect 43824 26450 43852 26862
rect 43812 26444 43864 26450
rect 43812 26386 43864 26392
rect 44744 26314 44772 28562
rect 45020 26382 45048 29242
rect 45836 28076 45888 28082
rect 45836 28018 45888 28024
rect 45284 27872 45336 27878
rect 45284 27814 45336 27820
rect 45296 26382 45324 27814
rect 45376 26920 45428 26926
rect 45376 26862 45428 26868
rect 45388 26586 45416 26862
rect 45744 26784 45796 26790
rect 45744 26726 45796 26732
rect 45376 26580 45428 26586
rect 45376 26522 45428 26528
rect 45560 26580 45612 26586
rect 45560 26522 45612 26528
rect 45008 26376 45060 26382
rect 45008 26318 45060 26324
rect 45284 26376 45336 26382
rect 45284 26318 45336 26324
rect 44732 26308 44784 26314
rect 44732 26250 44784 26256
rect 44272 25968 44324 25974
rect 44272 25910 44324 25916
rect 44284 25362 44312 25910
rect 44744 25838 44772 26250
rect 45020 25906 45048 26318
rect 45296 25906 45324 26318
rect 45008 25900 45060 25906
rect 45008 25842 45060 25848
rect 45284 25900 45336 25906
rect 45284 25842 45336 25848
rect 44732 25832 44784 25838
rect 44732 25774 44784 25780
rect 44364 25696 44416 25702
rect 44364 25638 44416 25644
rect 45376 25696 45428 25702
rect 45376 25638 45428 25644
rect 45468 25696 45520 25702
rect 45468 25638 45520 25644
rect 44376 25498 44404 25638
rect 44364 25492 44416 25498
rect 44364 25434 44416 25440
rect 44272 25356 44324 25362
rect 44272 25298 44324 25304
rect 44180 25288 44232 25294
rect 44180 25230 44232 25236
rect 43444 25220 43496 25226
rect 43444 25162 43496 25168
rect 44192 24818 44220 25230
rect 43260 24812 43312 24818
rect 43260 24754 43312 24760
rect 44180 24812 44232 24818
rect 44180 24754 44232 24760
rect 43272 23730 43300 24754
rect 44284 24698 44312 25298
rect 44376 24886 44404 25434
rect 45284 25424 45336 25430
rect 45284 25366 45336 25372
rect 44548 25356 44600 25362
rect 44548 25298 44600 25304
rect 44364 24880 44416 24886
rect 44364 24822 44416 24828
rect 44560 24818 44588 25298
rect 44916 25152 44968 25158
rect 44916 25094 44968 25100
rect 45192 25152 45244 25158
rect 45192 25094 45244 25100
rect 44548 24812 44600 24818
rect 44548 24754 44600 24760
rect 44364 24744 44416 24750
rect 44284 24692 44364 24698
rect 44284 24686 44416 24692
rect 44284 24670 44404 24686
rect 44732 24608 44784 24614
rect 44732 24550 44784 24556
rect 43904 24268 43956 24274
rect 43904 24210 43956 24216
rect 43812 24064 43864 24070
rect 43812 24006 43864 24012
rect 43168 23724 43220 23730
rect 43168 23666 43220 23672
rect 43260 23724 43312 23730
rect 43260 23666 43312 23672
rect 42800 23656 42852 23662
rect 42800 23598 42852 23604
rect 42536 22066 42656 22094
rect 42156 22024 42208 22030
rect 42156 21966 42208 21972
rect 42168 20534 42196 21966
rect 42156 20528 42208 20534
rect 42156 20470 42208 20476
rect 42064 19916 42116 19922
rect 42064 19858 42116 19864
rect 41880 19236 41932 19242
rect 41880 19178 41932 19184
rect 42064 19168 42116 19174
rect 42064 19110 42116 19116
rect 42076 18970 42104 19110
rect 42064 18964 42116 18970
rect 42064 18906 42116 18912
rect 42168 18850 42196 20470
rect 42340 19780 42392 19786
rect 42340 19722 42392 19728
rect 42352 18970 42380 19722
rect 42340 18964 42392 18970
rect 42340 18906 42392 18912
rect 41604 18828 41656 18834
rect 41604 18770 41656 18776
rect 42076 18822 42196 18850
rect 42076 18766 42104 18822
rect 42064 18760 42116 18766
rect 42064 18702 42116 18708
rect 42432 18216 42484 18222
rect 42432 18158 42484 18164
rect 42444 17814 42472 18158
rect 42432 17808 42484 17814
rect 42432 17750 42484 17756
rect 40500 17740 40552 17746
rect 40500 17682 40552 17688
rect 40960 17604 41012 17610
rect 40960 17546 41012 17552
rect 40408 17332 40460 17338
rect 40408 17274 40460 17280
rect 40972 17202 41000 17546
rect 41144 17536 41196 17542
rect 41144 17478 41196 17484
rect 41236 17536 41288 17542
rect 41236 17478 41288 17484
rect 41156 17202 41184 17478
rect 40960 17196 41012 17202
rect 40960 17138 41012 17144
rect 41144 17196 41196 17202
rect 41144 17138 41196 17144
rect 40224 17128 40276 17134
rect 40224 17070 40276 17076
rect 39856 16788 39908 16794
rect 39856 16730 39908 16736
rect 40236 16454 40264 17070
rect 40316 17060 40368 17066
rect 40316 17002 40368 17008
rect 40328 16574 40356 17002
rect 40972 16658 41000 17138
rect 41248 17066 41276 17478
rect 41236 17060 41288 17066
rect 41236 17002 41288 17008
rect 40960 16652 41012 16658
rect 40960 16594 41012 16600
rect 40408 16584 40460 16590
rect 40328 16546 40408 16574
rect 40408 16526 40460 16532
rect 40224 16448 40276 16454
rect 40224 16390 40276 16396
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 41420 11756 41472 11762
rect 41420 11698 41472 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 27160 9920 27212 9926
rect 27160 9862 27212 9868
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25516 3602 25544 3878
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 25596 3664 25648 3670
rect 25792 3618 25820 3674
rect 25648 3612 25820 3618
rect 25596 3606 25820 3612
rect 25504 3596 25556 3602
rect 25608 3590 25820 3606
rect 25504 3538 25556 3544
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 25332 3058 25360 3470
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 23860 800 23888 2382
rect 25792 800 25820 3402
rect 27172 2990 27200 9862
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 38660 4140 38712 4146
rect 38660 4082 38712 4088
rect 40776 4140 40828 4146
rect 40776 4082 40828 4088
rect 38568 4004 38620 4010
rect 38568 3946 38620 3952
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 28172 3664 28224 3670
rect 28356 3664 28408 3670
rect 28224 3612 28356 3618
rect 28172 3606 28408 3612
rect 28184 3590 28396 3606
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 27252 2984 27304 2990
rect 27252 2926 27304 2932
rect 27264 898 27292 2926
rect 27816 2582 27844 3470
rect 28356 3392 28408 3398
rect 28356 3334 28408 3340
rect 27804 2576 27856 2582
rect 27804 2518 27856 2524
rect 28368 2514 28396 3334
rect 32140 3058 32168 3470
rect 38476 3460 38528 3466
rect 38476 3402 38528 3408
rect 32312 3392 32364 3398
rect 32312 3334 32364 3340
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 32324 2990 32352 3334
rect 38488 3194 38516 3402
rect 38476 3188 38528 3194
rect 38476 3130 38528 3136
rect 38580 3058 38608 3946
rect 38568 3052 38620 3058
rect 38568 2994 38620 3000
rect 32312 2984 32364 2990
rect 32312 2926 32364 2932
rect 32404 2984 32456 2990
rect 32404 2926 32456 2932
rect 28356 2508 28408 2514
rect 28356 2450 28408 2456
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 26436 870 26648 898
rect 26436 800 26464 870
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 2566 0 2678 800
rect 3210 0 3322 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 11582 0 11694 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14158 0 14270 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 18022 0 18134 800
rect 19310 0 19422 800
rect 19954 0 20066 800
rect 20598 0 20710 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25750 0 25862 800
rect 26394 0 26506 800
rect 26620 762 26648 870
rect 26896 870 27292 898
rect 26896 762 26924 870
rect 27724 800 27752 2314
rect 32416 1578 32444 2926
rect 38672 2922 38700 4082
rect 38752 3936 38804 3942
rect 38752 3878 38804 3884
rect 40040 3936 40092 3942
rect 40040 3878 40092 3884
rect 38764 3126 38792 3878
rect 40052 3602 40080 3878
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 40592 3596 40644 3602
rect 40592 3538 40644 3544
rect 38752 3120 38804 3126
rect 38752 3062 38804 3068
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 38660 2916 38712 2922
rect 38660 2858 38712 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 32232 1550 32444 1578
rect 32232 800 32260 1550
rect 39316 800 39344 2926
rect 40604 800 40632 3538
rect 40788 3058 40816 4082
rect 41432 4010 41460 11698
rect 42340 4616 42392 4622
rect 42340 4558 42392 4564
rect 41512 4276 41564 4282
rect 41512 4218 41564 4224
rect 41524 4010 41552 4218
rect 41972 4208 42024 4214
rect 41972 4150 42024 4156
rect 41420 4004 41472 4010
rect 41420 3946 41472 3952
rect 41512 4004 41564 4010
rect 41512 3946 41564 3952
rect 40868 3936 40920 3942
rect 40868 3878 40920 3884
rect 41788 3936 41840 3942
rect 41788 3878 41840 3884
rect 40880 3126 40908 3878
rect 41800 3670 41828 3878
rect 41880 3732 41932 3738
rect 41880 3674 41932 3680
rect 41788 3664 41840 3670
rect 41788 3606 41840 3612
rect 40868 3120 40920 3126
rect 40868 3062 40920 3068
rect 40776 3052 40828 3058
rect 40776 2994 40828 3000
rect 41236 2916 41288 2922
rect 41236 2858 41288 2864
rect 41248 800 41276 2858
rect 41892 800 41920 3674
rect 41984 3602 42012 4150
rect 42156 3936 42208 3942
rect 42156 3878 42208 3884
rect 42168 3602 42196 3878
rect 41972 3596 42024 3602
rect 41972 3538 42024 3544
rect 42156 3596 42208 3602
rect 42156 3538 42208 3544
rect 42352 2514 42380 4558
rect 42536 4146 42564 22066
rect 42708 21956 42760 21962
rect 42708 21898 42760 21904
rect 42616 21888 42668 21894
rect 42616 21830 42668 21836
rect 42628 19718 42656 21830
rect 42720 21622 42748 21898
rect 42708 21616 42760 21622
rect 42708 21558 42760 21564
rect 42708 20800 42760 20806
rect 42812 20754 42840 23598
rect 43180 22094 43208 23666
rect 42996 22066 43208 22094
rect 42996 22030 43024 22066
rect 42984 22024 43036 22030
rect 42984 21966 43036 21972
rect 42984 21888 43036 21894
rect 42984 21830 43036 21836
rect 42996 21690 43024 21830
rect 42984 21684 43036 21690
rect 42984 21626 43036 21632
rect 42892 21548 42944 21554
rect 42892 21490 42944 21496
rect 42904 20806 42932 21490
rect 42996 20942 43024 21626
rect 43076 21548 43128 21554
rect 43076 21490 43128 21496
rect 43088 21146 43116 21490
rect 43076 21140 43128 21146
rect 43076 21082 43128 21088
rect 42984 20936 43036 20942
rect 42984 20878 43036 20884
rect 42760 20748 42840 20754
rect 42708 20742 42840 20748
rect 42892 20800 42944 20806
rect 42892 20742 42944 20748
rect 42720 20726 42840 20742
rect 42616 19712 42668 19718
rect 42616 19654 42668 19660
rect 42628 19378 42656 19654
rect 42616 19372 42668 19378
rect 42616 19314 42668 19320
rect 43180 18850 43208 22066
rect 43272 21350 43300 23666
rect 43824 23662 43852 24006
rect 43916 23730 43944 24210
rect 43996 24200 44048 24206
rect 43996 24142 44048 24148
rect 44008 23866 44036 24142
rect 44744 24138 44772 24550
rect 44732 24132 44784 24138
rect 44732 24074 44784 24080
rect 43996 23860 44048 23866
rect 43996 23802 44048 23808
rect 43904 23724 43956 23730
rect 43904 23666 43956 23672
rect 43812 23656 43864 23662
rect 43812 23598 43864 23604
rect 44180 22432 44232 22438
rect 44180 22374 44232 22380
rect 44192 22098 44220 22374
rect 44180 22092 44232 22098
rect 44180 22034 44232 22040
rect 44192 21554 44220 22034
rect 44548 22024 44600 22030
rect 44548 21966 44600 21972
rect 44272 21888 44324 21894
rect 44272 21830 44324 21836
rect 44180 21548 44232 21554
rect 44180 21490 44232 21496
rect 43260 21344 43312 21350
rect 43260 21286 43312 21292
rect 43260 19916 43312 19922
rect 43260 19858 43312 19864
rect 43272 19378 43300 19858
rect 43628 19712 43680 19718
rect 43628 19654 43680 19660
rect 43260 19372 43312 19378
rect 43260 19314 43312 19320
rect 43536 18964 43588 18970
rect 43536 18906 43588 18912
rect 42996 18822 43208 18850
rect 42616 18760 42668 18766
rect 42616 18702 42668 18708
rect 42628 18358 42656 18702
rect 42996 18358 43024 18822
rect 43076 18692 43128 18698
rect 43076 18634 43128 18640
rect 42616 18352 42668 18358
rect 42984 18352 43036 18358
rect 42668 18300 42748 18306
rect 42616 18294 42748 18300
rect 42984 18294 43036 18300
rect 42628 18278 42748 18294
rect 42720 17814 42748 18278
rect 42892 18080 42944 18086
rect 42892 18022 42944 18028
rect 42708 17808 42760 17814
rect 42708 17750 42760 17756
rect 42720 17134 42748 17750
rect 42904 17746 42932 18022
rect 43088 17814 43116 18634
rect 43168 18624 43220 18630
rect 43168 18566 43220 18572
rect 43076 17808 43128 17814
rect 43076 17750 43128 17756
rect 43180 17746 43208 18566
rect 43548 18290 43576 18906
rect 43640 18834 43668 19654
rect 43628 18828 43680 18834
rect 43628 18770 43680 18776
rect 43536 18284 43588 18290
rect 43536 18226 43588 18232
rect 42892 17740 42944 17746
rect 42892 17682 42944 17688
rect 43168 17740 43220 17746
rect 43168 17682 43220 17688
rect 42984 17672 43036 17678
rect 42984 17614 43036 17620
rect 42996 17134 43024 17614
rect 43640 17202 43668 18770
rect 44284 18766 44312 21830
rect 44560 21622 44588 21966
rect 44732 21956 44784 21962
rect 44732 21898 44784 21904
rect 44744 21622 44772 21898
rect 44928 21690 44956 25094
rect 45100 24064 45152 24070
rect 45100 24006 45152 24012
rect 45008 23588 45060 23594
rect 45008 23530 45060 23536
rect 45020 23118 45048 23530
rect 45008 23112 45060 23118
rect 45008 23054 45060 23060
rect 45112 22710 45140 24006
rect 45100 22704 45152 22710
rect 45100 22646 45152 22652
rect 45008 22636 45060 22642
rect 45008 22578 45060 22584
rect 45020 22098 45048 22578
rect 45008 22092 45060 22098
rect 45008 22034 45060 22040
rect 44916 21684 44968 21690
rect 44916 21626 44968 21632
rect 44548 21616 44600 21622
rect 44548 21558 44600 21564
rect 44732 21616 44784 21622
rect 44732 21558 44784 21564
rect 44560 21486 44588 21558
rect 44364 21480 44416 21486
rect 44364 21422 44416 21428
rect 44548 21480 44600 21486
rect 44548 21422 44600 21428
rect 44376 21078 44404 21422
rect 44364 21072 44416 21078
rect 44364 21014 44416 21020
rect 44744 21010 44772 21558
rect 44916 21548 44968 21554
rect 44916 21490 44968 21496
rect 44824 21072 44876 21078
rect 44824 21014 44876 21020
rect 44732 21004 44784 21010
rect 44732 20946 44784 20952
rect 44744 20398 44772 20946
rect 44836 20466 44864 21014
rect 44928 20466 44956 21490
rect 45020 21350 45048 22034
rect 45100 21480 45152 21486
rect 45100 21422 45152 21428
rect 45008 21344 45060 21350
rect 45008 21286 45060 21292
rect 45020 20942 45048 21286
rect 45112 21146 45140 21422
rect 45204 21146 45232 25094
rect 45296 24818 45324 25366
rect 45388 25294 45416 25638
rect 45480 25430 45508 25638
rect 45468 25424 45520 25430
rect 45468 25366 45520 25372
rect 45376 25288 45428 25294
rect 45428 25248 45508 25276
rect 45376 25230 45428 25236
rect 45480 24818 45508 25248
rect 45572 25226 45600 26522
rect 45652 26444 45704 26450
rect 45652 26386 45704 26392
rect 45560 25220 45612 25226
rect 45560 25162 45612 25168
rect 45572 24886 45600 25162
rect 45560 24880 45612 24886
rect 45560 24822 45612 24828
rect 45284 24812 45336 24818
rect 45284 24754 45336 24760
rect 45468 24812 45520 24818
rect 45468 24754 45520 24760
rect 45560 24676 45612 24682
rect 45560 24618 45612 24624
rect 45468 24608 45520 24614
rect 45468 24550 45520 24556
rect 45480 24206 45508 24550
rect 45468 24200 45520 24206
rect 45468 24142 45520 24148
rect 45572 23905 45600 24618
rect 45558 23896 45614 23905
rect 45558 23831 45614 23840
rect 45664 23118 45692 26386
rect 45756 26382 45784 26726
rect 45848 26518 45876 28018
rect 45940 26586 45968 31726
rect 46124 31414 46152 32710
rect 46480 32292 46532 32298
rect 46480 32234 46532 32240
rect 46492 31890 46520 32234
rect 46480 31884 46532 31890
rect 46480 31826 46532 31832
rect 46676 31754 46704 36518
rect 46756 36236 46808 36242
rect 46756 36178 46808 36184
rect 46768 35154 46796 36178
rect 46860 36174 46888 36518
rect 46952 36378 46980 37606
rect 47032 36780 47084 36786
rect 47032 36722 47084 36728
rect 46940 36372 46992 36378
rect 46940 36314 46992 36320
rect 46848 36168 46900 36174
rect 46848 36110 46900 36116
rect 46952 35698 46980 36314
rect 47044 35834 47072 36722
rect 47032 35828 47084 35834
rect 47032 35770 47084 35776
rect 46940 35692 46992 35698
rect 46940 35634 46992 35640
rect 46756 35148 46808 35154
rect 46756 35090 46808 35096
rect 46768 34066 46796 35090
rect 46848 35080 46900 35086
rect 46848 35022 46900 35028
rect 46860 34746 46888 35022
rect 46848 34740 46900 34746
rect 46848 34682 46900 34688
rect 46756 34060 46808 34066
rect 46756 34002 46808 34008
rect 46848 33516 46900 33522
rect 46848 33458 46900 33464
rect 46860 33425 46888 33458
rect 46846 33416 46902 33425
rect 46846 33351 46902 33360
rect 46940 33312 46992 33318
rect 46940 33254 46992 33260
rect 46952 31958 46980 33254
rect 46940 31952 46992 31958
rect 46940 31894 46992 31900
rect 46584 31726 46704 31754
rect 46112 31408 46164 31414
rect 46112 31350 46164 31356
rect 46020 31340 46072 31346
rect 46020 31282 46072 31288
rect 46032 30938 46060 31282
rect 46020 30932 46072 30938
rect 46020 30874 46072 30880
rect 46124 30734 46152 31350
rect 46112 30728 46164 30734
rect 46112 30670 46164 30676
rect 46296 29640 46348 29646
rect 46296 29582 46348 29588
rect 46308 29170 46336 29582
rect 46480 29572 46532 29578
rect 46480 29514 46532 29520
rect 46296 29164 46348 29170
rect 46296 29106 46348 29112
rect 46492 28218 46520 29514
rect 46480 28212 46532 28218
rect 46480 28154 46532 28160
rect 46388 28076 46440 28082
rect 46388 28018 46440 28024
rect 46020 27396 46072 27402
rect 46020 27338 46072 27344
rect 45928 26580 45980 26586
rect 45928 26522 45980 26528
rect 45836 26512 45888 26518
rect 46032 26466 46060 27338
rect 46112 26988 46164 26994
rect 46112 26930 46164 26936
rect 45836 26454 45888 26460
rect 45940 26438 46060 26466
rect 45940 26382 45968 26438
rect 45744 26376 45796 26382
rect 45744 26318 45796 26324
rect 45928 26376 45980 26382
rect 45928 26318 45980 26324
rect 45756 25906 45784 26318
rect 45744 25900 45796 25906
rect 45744 25842 45796 25848
rect 45836 24608 45888 24614
rect 45836 24550 45888 24556
rect 45848 23730 45876 24550
rect 45836 23724 45888 23730
rect 45836 23666 45888 23672
rect 45284 23112 45336 23118
rect 45284 23054 45336 23060
rect 45652 23112 45704 23118
rect 45652 23054 45704 23060
rect 45296 21894 45324 23054
rect 45376 22704 45428 22710
rect 45376 22646 45428 22652
rect 45388 22030 45416 22646
rect 45652 22432 45704 22438
rect 45652 22374 45704 22380
rect 45376 22024 45428 22030
rect 45376 21966 45428 21972
rect 45468 22024 45520 22030
rect 45468 21966 45520 21972
rect 45284 21888 45336 21894
rect 45284 21830 45336 21836
rect 45284 21684 45336 21690
rect 45284 21626 45336 21632
rect 45100 21140 45152 21146
rect 45100 21082 45152 21088
rect 45192 21140 45244 21146
rect 45192 21082 45244 21088
rect 45008 20936 45060 20942
rect 45008 20878 45060 20884
rect 44824 20460 44876 20466
rect 44824 20402 44876 20408
rect 44916 20460 44968 20466
rect 44916 20402 44968 20408
rect 44732 20392 44784 20398
rect 44732 20334 44784 20340
rect 44456 19916 44508 19922
rect 44456 19858 44508 19864
rect 44364 19712 44416 19718
rect 44364 19654 44416 19660
rect 44376 18902 44404 19654
rect 44364 18896 44416 18902
rect 44364 18838 44416 18844
rect 44272 18760 44324 18766
rect 44272 18702 44324 18708
rect 44088 18692 44140 18698
rect 44088 18634 44140 18640
rect 44100 18154 44128 18634
rect 44180 18352 44232 18358
rect 44180 18294 44232 18300
rect 44088 18148 44140 18154
rect 44088 18090 44140 18096
rect 44100 17610 44128 18090
rect 44088 17604 44140 17610
rect 44088 17546 44140 17552
rect 44100 17202 44128 17546
rect 44192 17338 44220 18294
rect 44284 17678 44312 18702
rect 44468 18426 44496 19858
rect 44836 19854 44864 20402
rect 45296 19854 45324 21626
rect 45388 20942 45416 21966
rect 45376 20936 45428 20942
rect 45376 20878 45428 20884
rect 45480 20602 45508 21966
rect 45560 21888 45612 21894
rect 45560 21830 45612 21836
rect 45468 20596 45520 20602
rect 45468 20538 45520 20544
rect 45572 20534 45600 21830
rect 45664 21554 45692 22374
rect 45940 22094 45968 26318
rect 46124 24188 46152 26930
rect 46296 26784 46348 26790
rect 46296 26726 46348 26732
rect 46202 26616 46258 26625
rect 46202 26551 46258 26560
rect 46216 24342 46244 26551
rect 46308 26450 46336 26726
rect 46296 26444 46348 26450
rect 46296 26386 46348 26392
rect 46204 24336 46256 24342
rect 46204 24278 46256 24284
rect 46124 24160 46244 24188
rect 46020 23724 46072 23730
rect 46020 23666 46072 23672
rect 46112 23724 46164 23730
rect 46112 23666 46164 23672
rect 45848 22066 45968 22094
rect 45652 21548 45704 21554
rect 45652 21490 45704 21496
rect 45560 20528 45612 20534
rect 45480 20476 45560 20482
rect 45480 20470 45612 20476
rect 45480 20454 45600 20470
rect 45480 20058 45508 20454
rect 45572 20405 45600 20454
rect 45468 20052 45520 20058
rect 45468 19994 45520 20000
rect 44824 19848 44876 19854
rect 44824 19790 44876 19796
rect 45284 19848 45336 19854
rect 45284 19790 45336 19796
rect 45192 19780 45244 19786
rect 45192 19722 45244 19728
rect 45204 19378 45232 19722
rect 44640 19372 44692 19378
rect 44640 19314 44692 19320
rect 45008 19372 45060 19378
rect 45008 19314 45060 19320
rect 45192 19372 45244 19378
rect 45192 19314 45244 19320
rect 44652 18970 44680 19314
rect 44640 18964 44692 18970
rect 44640 18906 44692 18912
rect 44732 18624 44784 18630
rect 44732 18566 44784 18572
rect 44456 18420 44508 18426
rect 44456 18362 44508 18368
rect 44744 18290 44772 18566
rect 45020 18426 45048 19314
rect 45468 18896 45520 18902
rect 45468 18838 45520 18844
rect 45008 18420 45060 18426
rect 45008 18362 45060 18368
rect 44732 18284 44784 18290
rect 44732 18226 44784 18232
rect 45480 18222 45508 18838
rect 45468 18216 45520 18222
rect 45468 18158 45520 18164
rect 45560 17876 45612 17882
rect 45560 17818 45612 17824
rect 45572 17785 45600 17818
rect 45558 17776 45614 17785
rect 45558 17711 45614 17720
rect 44272 17672 44324 17678
rect 44272 17614 44324 17620
rect 44180 17332 44232 17338
rect 44180 17274 44232 17280
rect 44284 17202 44312 17614
rect 43628 17196 43680 17202
rect 43628 17138 43680 17144
rect 44088 17196 44140 17202
rect 44088 17138 44140 17144
rect 44272 17196 44324 17202
rect 44272 17138 44324 17144
rect 42708 17128 42760 17134
rect 42708 17070 42760 17076
rect 42984 17128 43036 17134
rect 42984 17070 43036 17076
rect 45848 8634 45876 22066
rect 46032 20942 46060 23666
rect 46124 23322 46152 23666
rect 46112 23316 46164 23322
rect 46112 23258 46164 23264
rect 46112 21344 46164 21350
rect 46112 21286 46164 21292
rect 46124 20942 46152 21286
rect 46020 20936 46072 20942
rect 45940 20896 46020 20924
rect 45940 19174 45968 20896
rect 46020 20878 46072 20884
rect 46112 20936 46164 20942
rect 46112 20878 46164 20884
rect 46020 19508 46072 19514
rect 46020 19450 46072 19456
rect 45928 19168 45980 19174
rect 45928 19110 45980 19116
rect 46032 18834 46060 19450
rect 46020 18828 46072 18834
rect 46020 18770 46072 18776
rect 46032 18290 46060 18770
rect 46020 18284 46072 18290
rect 46020 18226 46072 18232
rect 45836 8628 45888 8634
rect 45836 8570 45888 8576
rect 45560 6316 45612 6322
rect 45560 6258 45612 6264
rect 45376 4480 45428 4486
rect 45376 4422 45428 4428
rect 45388 4214 45416 4422
rect 45572 4282 45600 6258
rect 45652 5704 45704 5710
rect 45652 5646 45704 5652
rect 45836 5704 45888 5710
rect 45836 5646 45888 5652
rect 45560 4276 45612 4282
rect 45560 4218 45612 4224
rect 45376 4208 45428 4214
rect 45376 4150 45428 4156
rect 42524 4140 42576 4146
rect 42524 4082 42576 4088
rect 43628 3936 43680 3942
rect 43628 3878 43680 3884
rect 44732 3936 44784 3942
rect 44732 3878 44784 3884
rect 43352 3460 43404 3466
rect 43352 3402 43404 3408
rect 43364 2922 43392 3402
rect 43640 2990 43668 3878
rect 44744 3058 44772 3878
rect 45664 3738 45692 5646
rect 45848 4826 45876 5646
rect 45836 4820 45888 4826
rect 45836 4762 45888 4768
rect 46216 4622 46244 24160
rect 46296 23724 46348 23730
rect 46296 23666 46348 23672
rect 46308 20942 46336 23666
rect 46296 20936 46348 20942
rect 46296 20878 46348 20884
rect 46308 19718 46336 20878
rect 46296 19712 46348 19718
rect 46296 19654 46348 19660
rect 46296 18760 46348 18766
rect 46296 18702 46348 18708
rect 46308 18358 46336 18702
rect 46296 18352 46348 18358
rect 46296 18294 46348 18300
rect 46296 6112 46348 6118
rect 46296 6054 46348 6060
rect 46308 5302 46336 6054
rect 46296 5296 46348 5302
rect 46296 5238 46348 5244
rect 46296 5024 46348 5030
rect 46296 4966 46348 4972
rect 46308 4690 46336 4966
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 46204 4616 46256 4622
rect 46204 4558 46256 4564
rect 45652 3732 45704 3738
rect 45652 3674 45704 3680
rect 46400 3670 46428 28018
rect 46480 27872 46532 27878
rect 46480 27814 46532 27820
rect 46492 27538 46520 27814
rect 46480 27532 46532 27538
rect 46480 27474 46532 27480
rect 46480 25696 46532 25702
rect 46480 25638 46532 25644
rect 46492 25362 46520 25638
rect 46480 25356 46532 25362
rect 46480 25298 46532 25304
rect 46584 20466 46612 31726
rect 46940 31680 46992 31686
rect 46940 31622 46992 31628
rect 46848 31340 46900 31346
rect 46952 31328 46980 31622
rect 47032 31408 47084 31414
rect 47032 31350 47084 31356
rect 46900 31300 46980 31328
rect 46848 31282 46900 31288
rect 47044 30938 47072 31350
rect 47032 30932 47084 30938
rect 47032 30874 47084 30880
rect 47044 30394 47072 30874
rect 47032 30388 47084 30394
rect 47032 30330 47084 30336
rect 46846 29336 46902 29345
rect 46846 29271 46902 29280
rect 46860 27538 46888 29271
rect 46940 28484 46992 28490
rect 46940 28426 46992 28432
rect 46848 27532 46900 27538
rect 46848 27474 46900 27480
rect 46952 27130 46980 28426
rect 46940 27124 46992 27130
rect 46940 27066 46992 27072
rect 46940 26512 46992 26518
rect 46940 26454 46992 26460
rect 46952 25906 46980 26454
rect 46940 25900 46992 25906
rect 46940 25842 46992 25848
rect 46756 25356 46808 25362
rect 46756 25298 46808 25304
rect 46664 23112 46716 23118
rect 46664 23054 46716 23060
rect 46676 21026 46704 23054
rect 46768 21865 46796 25298
rect 47032 24812 47084 24818
rect 47032 24754 47084 24760
rect 46940 24132 46992 24138
rect 46940 24074 46992 24080
rect 46952 23866 46980 24074
rect 46940 23860 46992 23866
rect 46940 23802 46992 23808
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 46952 23118 46980 23462
rect 47044 23322 47072 24754
rect 47032 23316 47084 23322
rect 47032 23258 47084 23264
rect 46940 23112 46992 23118
rect 46940 23054 46992 23060
rect 47032 22432 47084 22438
rect 47032 22374 47084 22380
rect 47044 22098 47072 22374
rect 47032 22092 47084 22098
rect 47032 22034 47084 22040
rect 46754 21856 46810 21865
rect 46754 21791 46810 21800
rect 46676 21010 46796 21026
rect 46676 21004 46808 21010
rect 46676 20998 46756 21004
rect 46756 20946 46808 20952
rect 46572 20460 46624 20466
rect 46572 20402 46624 20408
rect 46480 20256 46532 20262
rect 46480 20198 46532 20204
rect 46492 19922 46520 20198
rect 46480 19916 46532 19922
rect 46480 19858 46532 19864
rect 46768 19378 46796 20946
rect 46756 19372 46808 19378
rect 46756 19314 46808 19320
rect 46940 18692 46992 18698
rect 46940 18634 46992 18640
rect 46952 18426 46980 18634
rect 46940 18420 46992 18426
rect 46940 18362 46992 18368
rect 46940 16992 46992 16998
rect 46940 16934 46992 16940
rect 46952 16522 46980 16934
rect 46940 16516 46992 16522
rect 46940 16458 46992 16464
rect 46480 14816 46532 14822
rect 46480 14758 46532 14764
rect 46492 14482 46520 14758
rect 46480 14476 46532 14482
rect 46480 14418 46532 14424
rect 47136 13802 47164 45766
rect 47228 23730 47256 46106
rect 47676 45892 47728 45898
rect 47676 45834 47728 45840
rect 47688 45558 47716 45834
rect 47676 45552 47728 45558
rect 47676 45494 47728 45500
rect 47308 45484 47360 45490
rect 47308 45426 47360 45432
rect 47320 38434 47348 45426
rect 47584 44736 47636 44742
rect 47584 44678 47636 44684
rect 47596 43314 47624 44678
rect 47860 44396 47912 44402
rect 47860 44338 47912 44344
rect 47584 43308 47636 43314
rect 47584 43250 47636 43256
rect 47596 38962 47624 43250
rect 47676 43104 47728 43110
rect 47676 43046 47728 43052
rect 47688 42770 47716 43046
rect 47676 42764 47728 42770
rect 47676 42706 47728 42712
rect 47768 39840 47820 39846
rect 47768 39782 47820 39788
rect 47780 39506 47808 39782
rect 47768 39500 47820 39506
rect 47768 39442 47820 39448
rect 47676 39364 47728 39370
rect 47676 39306 47728 39312
rect 47688 39098 47716 39306
rect 47676 39092 47728 39098
rect 47676 39034 47728 39040
rect 47584 38956 47636 38962
rect 47584 38898 47636 38904
rect 47320 38406 47624 38434
rect 47400 38344 47452 38350
rect 47398 38312 47400 38321
rect 47452 38312 47454 38321
rect 47398 38247 47454 38256
rect 47308 32836 47360 32842
rect 47308 32778 47360 32784
rect 47320 31346 47348 32778
rect 47308 31340 47360 31346
rect 47308 31282 47360 31288
rect 47216 23724 47268 23730
rect 47216 23666 47268 23672
rect 47412 17202 47440 38247
rect 47492 38208 47544 38214
rect 47492 38150 47544 38156
rect 47504 37194 47532 38150
rect 47492 37188 47544 37194
rect 47492 37130 47544 37136
rect 47596 32994 47624 38406
rect 47768 35692 47820 35698
rect 47768 35634 47820 35640
rect 47780 34678 47808 35634
rect 47768 34672 47820 34678
rect 47768 34614 47820 34620
rect 47676 33924 47728 33930
rect 47676 33866 47728 33872
rect 47688 33114 47716 33866
rect 47676 33108 47728 33114
rect 47676 33050 47728 33056
rect 47596 32966 47716 32994
rect 47584 32224 47636 32230
rect 47584 32166 47636 32172
rect 47492 31476 47544 31482
rect 47492 31418 47544 31424
rect 47504 30938 47532 31418
rect 47492 30932 47544 30938
rect 47492 30874 47544 30880
rect 47596 30734 47624 32166
rect 47584 30728 47636 30734
rect 47584 30670 47636 30676
rect 47688 28778 47716 32966
rect 47768 32428 47820 32434
rect 47768 32370 47820 32376
rect 47780 31482 47808 32370
rect 47768 31476 47820 31482
rect 47768 31418 47820 31424
rect 47768 31204 47820 31210
rect 47768 31146 47820 31152
rect 47780 30258 47808 31146
rect 47768 30252 47820 30258
rect 47768 30194 47820 30200
rect 47596 28750 47716 28778
rect 47596 26994 47624 28750
rect 47676 28620 47728 28626
rect 47676 28562 47728 28568
rect 47688 26994 47716 28562
rect 47768 27872 47820 27878
rect 47768 27814 47820 27820
rect 47780 27606 47808 27814
rect 47768 27600 47820 27606
rect 47768 27542 47820 27548
rect 47584 26988 47636 26994
rect 47584 26930 47636 26936
rect 47676 26988 47728 26994
rect 47676 26930 47728 26936
rect 47768 25220 47820 25226
rect 47768 25162 47820 25168
rect 47780 24818 47808 25162
rect 47768 24812 47820 24818
rect 47768 24754 47820 24760
rect 47768 24268 47820 24274
rect 47768 24210 47820 24216
rect 47780 23730 47808 24210
rect 47768 23724 47820 23730
rect 47768 23666 47820 23672
rect 47676 22432 47728 22438
rect 47676 22374 47728 22380
rect 47688 21962 47716 22374
rect 47676 21956 47728 21962
rect 47676 21898 47728 21904
rect 47676 21480 47728 21486
rect 47676 21422 47728 21428
rect 47688 21146 47716 21422
rect 47676 21140 47728 21146
rect 47676 21082 47728 21088
rect 47768 19780 47820 19786
rect 47768 19722 47820 19728
rect 47780 19310 47808 19722
rect 47768 19304 47820 19310
rect 47768 19246 47820 19252
rect 47872 18222 47900 44338
rect 48056 43858 48084 49286
rect 48290 49200 48402 50000
rect 48934 49200 49046 50000
rect 49578 49200 49690 50000
rect 48332 46034 48360 49200
rect 48320 46028 48372 46034
rect 48320 45970 48372 45976
rect 48134 44976 48190 44985
rect 48134 44911 48136 44920
rect 48188 44911 48190 44920
rect 48136 44882 48188 44888
rect 48044 43852 48096 43858
rect 48044 43794 48096 43800
rect 48136 42628 48188 42634
rect 48136 42570 48188 42576
rect 48148 41585 48176 42570
rect 48134 41576 48190 41585
rect 48134 41511 48190 41520
rect 48228 41540 48280 41546
rect 48228 41482 48280 41488
rect 48136 40452 48188 40458
rect 48136 40394 48188 40400
rect 48148 39545 48176 40394
rect 48134 39536 48190 39545
rect 48134 39471 48190 39480
rect 48136 39364 48188 39370
rect 48136 39306 48188 39312
rect 48148 38185 48176 39306
rect 48134 38176 48190 38185
rect 48134 38111 48190 38120
rect 48240 37505 48268 41482
rect 48226 37496 48282 37505
rect 48226 37431 48282 37440
rect 48136 37188 48188 37194
rect 48136 37130 48188 37136
rect 48148 36145 48176 37130
rect 48134 36136 48190 36145
rect 48134 36071 48190 36080
rect 48044 33856 48096 33862
rect 48044 33798 48096 33804
rect 48056 31686 48084 33798
rect 48134 32736 48190 32745
rect 48134 32671 48190 32680
rect 48148 31890 48176 32671
rect 48136 31884 48188 31890
rect 48136 31826 48188 31832
rect 48044 31680 48096 31686
rect 48044 31622 48096 31628
rect 48056 31278 48084 31622
rect 48044 31272 48096 31278
rect 48044 31214 48096 31220
rect 48136 29572 48188 29578
rect 48136 29514 48188 29520
rect 48148 28665 48176 29514
rect 48134 28656 48190 28665
rect 48134 28591 48190 28600
rect 48136 28484 48188 28490
rect 48136 28426 48188 28432
rect 48148 27985 48176 28426
rect 48134 27976 48190 27985
rect 48134 27911 48190 27920
rect 48134 25936 48190 25945
rect 48134 25871 48190 25880
rect 48148 24274 48176 25871
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 48134 22536 48190 22545
rect 48134 22471 48190 22480
rect 48148 22098 48176 22471
rect 48136 22092 48188 22098
rect 48136 22034 48188 22040
rect 48136 21548 48188 21554
rect 48136 21490 48188 21496
rect 48148 21146 48176 21490
rect 48136 21140 48188 21146
rect 48136 21082 48188 21088
rect 48134 20496 48190 20505
rect 48134 20431 48190 20440
rect 48148 19922 48176 20431
rect 48136 19916 48188 19922
rect 48136 19858 48188 19864
rect 48134 19136 48190 19145
rect 48134 19071 48190 19080
rect 48148 18834 48176 19071
rect 48136 18828 48188 18834
rect 48136 18770 48188 18776
rect 47860 18216 47912 18222
rect 47860 18158 47912 18164
rect 47400 17196 47452 17202
rect 47400 17138 47452 17144
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 47768 16992 47820 16998
rect 47768 16934 47820 16940
rect 47780 16658 47808 16934
rect 48148 16658 48176 17031
rect 47768 16652 47820 16658
rect 47768 16594 47820 16600
rect 48136 16652 48188 16658
rect 48136 16594 48188 16600
rect 47676 15496 47728 15502
rect 47676 15438 47728 15444
rect 47584 15020 47636 15026
rect 47584 14962 47636 14968
rect 46664 13796 46716 13802
rect 46664 13738 46716 13744
rect 47124 13796 47176 13802
rect 47124 13738 47176 13744
rect 46676 12850 46704 13738
rect 47596 12850 47624 14962
rect 47688 14550 47716 15438
rect 48134 15056 48190 15065
rect 48134 14991 48190 15000
rect 47676 14544 47728 14550
rect 47676 14486 47728 14492
rect 48148 14482 48176 14991
rect 48136 14476 48188 14482
rect 48136 14418 48188 14424
rect 47768 13728 47820 13734
rect 47768 13670 47820 13676
rect 48134 13696 48190 13705
rect 47780 13394 47808 13670
rect 48134 13631 48190 13640
rect 48148 13394 48176 13631
rect 47768 13388 47820 13394
rect 47768 13330 47820 13336
rect 48136 13388 48188 13394
rect 48136 13330 48188 13336
rect 47676 13252 47728 13258
rect 47676 13194 47728 13200
rect 47688 12986 47716 13194
rect 48134 13016 48190 13025
rect 47676 12980 47728 12986
rect 48134 12951 48190 12960
rect 47676 12922 47728 12928
rect 46664 12844 46716 12850
rect 46664 12786 46716 12792
rect 47584 12844 47636 12850
rect 47584 12786 47636 12792
rect 46480 12640 46532 12646
rect 46480 12582 46532 12588
rect 46492 12306 46520 12582
rect 46480 12300 46532 12306
rect 46480 12242 46532 12248
rect 46480 11552 46532 11558
rect 46480 11494 46532 11500
rect 46492 11218 46520 11494
rect 46480 11212 46532 11218
rect 46480 11154 46532 11160
rect 46676 6322 46704 12786
rect 47032 12640 47084 12646
rect 47032 12582 47084 12588
rect 47044 12374 47072 12582
rect 47596 12434 47624 12786
rect 47504 12406 47624 12434
rect 47032 12368 47084 12374
rect 46846 12336 46902 12345
rect 47032 12310 47084 12316
rect 46846 12271 46902 12280
rect 46860 11218 46888 12271
rect 46848 11212 46900 11218
rect 46848 11154 46900 11160
rect 47504 6390 47532 12406
rect 48148 12306 48176 12951
rect 48136 12300 48188 12306
rect 48136 12242 48188 12248
rect 47768 11552 47820 11558
rect 47768 11494 47820 11500
rect 47780 11286 47808 11494
rect 47768 11280 47820 11286
rect 47768 11222 47820 11228
rect 47952 8492 48004 8498
rect 47952 8434 48004 8440
rect 47964 8265 47992 8434
rect 47950 8256 48006 8265
rect 47950 8191 48006 8200
rect 47584 7404 47636 7410
rect 47584 7346 47636 7352
rect 47492 6384 47544 6390
rect 47492 6326 47544 6332
rect 46664 6316 46716 6322
rect 46664 6258 46716 6264
rect 46940 6112 46992 6118
rect 46940 6054 46992 6060
rect 46848 5160 46900 5166
rect 46848 5102 46900 5108
rect 46388 3664 46440 3670
rect 46388 3606 46440 3612
rect 45836 3528 45888 3534
rect 45836 3470 45888 3476
rect 45192 3392 45244 3398
rect 45192 3334 45244 3340
rect 44732 3052 44784 3058
rect 44732 2994 44784 3000
rect 43628 2984 43680 2990
rect 43628 2926 43680 2932
rect 43352 2916 43404 2922
rect 43352 2858 43404 2864
rect 42616 2848 42668 2854
rect 42616 2790 42668 2796
rect 42628 2514 42656 2790
rect 45204 2514 45232 3334
rect 45744 2916 45796 2922
rect 45744 2858 45796 2864
rect 42340 2508 42392 2514
rect 42340 2450 42392 2456
rect 42616 2508 42668 2514
rect 42616 2450 42668 2456
rect 45192 2508 45244 2514
rect 45192 2450 45244 2456
rect 45284 2508 45336 2514
rect 45284 2450 45336 2456
rect 45296 1306 45324 2450
rect 45112 1278 45324 1306
rect 45112 800 45140 1278
rect 45756 800 45784 2858
rect 45848 2582 45876 3470
rect 46572 2984 46624 2990
rect 46572 2926 46624 2932
rect 45836 2576 45888 2582
rect 45836 2518 45888 2524
rect 26620 734 26924 762
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 28970 0 29082 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 34122 0 34234 800
rect 34766 0 34878 800
rect 35410 0 35522 800
rect 36698 0 36810 800
rect 37342 0 37454 800
rect 38630 0 38742 800
rect 39274 0 39386 800
rect 40562 0 40674 800
rect 41206 0 41318 800
rect 41850 0 41962 800
rect 43138 0 43250 800
rect 43782 0 43894 800
rect 45070 0 45182 800
rect 45714 0 45826 800
rect 46584 105 46612 2926
rect 46860 2145 46888 5102
rect 46952 4690 46980 6054
rect 46940 4684 46992 4690
rect 46940 4626 46992 4632
rect 47032 4072 47084 4078
rect 47032 4014 47084 4020
rect 46846 2136 46902 2145
rect 46846 2071 46902 2080
rect 47044 800 47072 4014
rect 47596 3942 47624 7346
rect 47676 7200 47728 7206
rect 47676 7142 47728 7148
rect 47688 6866 47716 7142
rect 48134 6896 48190 6905
rect 47676 6860 47728 6866
rect 48134 6831 48136 6840
rect 47676 6802 47728 6808
rect 48188 6831 48190 6840
rect 48136 6802 48188 6808
rect 47768 6724 47820 6730
rect 47768 6666 47820 6672
rect 47780 6322 47808 6666
rect 47768 6316 47820 6322
rect 47768 6258 47820 6264
rect 48228 5636 48280 5642
rect 48228 5578 48280 5584
rect 48134 5536 48190 5545
rect 48134 5471 48190 5480
rect 48148 4690 48176 5471
rect 48136 4684 48188 4690
rect 48136 4626 48188 4632
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 47492 3596 47544 3602
rect 47492 3538 47544 3544
rect 47768 3596 47820 3602
rect 47768 3538 47820 3544
rect 47504 2650 47532 3538
rect 47676 3460 47728 3466
rect 47676 3402 47728 3408
rect 47688 3194 47716 3402
rect 47676 3188 47728 3194
rect 47676 3130 47728 3136
rect 47492 2644 47544 2650
rect 47492 2586 47544 2592
rect 47780 1714 47808 3538
rect 47688 1686 47808 1714
rect 47688 800 47716 1686
rect 48240 1465 48268 5578
rect 48964 2372 49016 2378
rect 48964 2314 49016 2320
rect 48226 1456 48282 1465
rect 48226 1391 48282 1400
rect 48976 800 49004 2314
rect 46570 96 46626 105
rect 46570 31 46626 40
rect 47002 0 47114 800
rect 47646 0 47758 800
rect 48934 0 49046 800
rect 49578 0 49690 800
<< via2 >>
rect 3606 48320 3662 48376
rect 2778 47640 2834 47696
rect 1674 46280 1730 46336
rect 2778 32680 2834 32736
rect 3330 41520 3386 41576
rect 3422 40840 3478 40896
rect 2778 25200 2834 25256
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3698 45600 3754 45656
rect 2778 23840 2834 23896
rect 2778 21800 2834 21856
rect 2778 20440 2834 20496
rect 2778 18400 2834 18456
rect 2778 17076 2780 17096
rect 2780 17076 2832 17096
rect 2832 17076 2834 17096
rect 2778 17040 2834 17076
rect 2778 15000 2834 15056
rect 2778 14320 2834 14376
rect 2778 11636 2780 11656
rect 2780 11636 2832 11656
rect 2832 11636 2834 11656
rect 2778 11600 2834 11636
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 3974 43560 4030 43616
rect 3238 10240 3294 10296
rect 2870 9560 2926 9616
rect 2778 7520 2834 7576
rect 2778 6840 2834 6896
rect 2870 5480 2926 5536
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3146 4800 3202 4856
rect 1858 3440 1914 3496
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 2760 4122 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 2778 1400 2834 1456
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 24122 27396 24178 27432
rect 24122 27376 24124 27396
rect 24124 27376 24176 27396
rect 24176 27376 24178 27396
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 33874 40996 33930 41032
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 33874 40976 33876 40996
rect 33876 40976 33928 40996
rect 33928 40976 33930 40996
rect 34794 40976 34850 41032
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 25594 29588 25596 29608
rect 25596 29588 25648 29608
rect 25648 29588 25650 29608
rect 25594 29552 25650 29588
rect 25778 29044 25780 29064
rect 25780 29044 25832 29064
rect 25832 29044 25834 29064
rect 25778 29008 25834 29044
rect 26146 29008 26202 29064
rect 28078 29552 28134 29608
rect 26514 27376 26570 27432
rect 32310 33088 32366 33144
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 33138 33108 33194 33144
rect 33138 33088 33140 33108
rect 33140 33088 33192 33108
rect 33192 33088 33194 33108
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 31942 28092 31944 28112
rect 31944 28092 31996 28112
rect 31996 28092 31998 28112
rect 31942 28056 31998 28092
rect 30562 27376 30618 27432
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 36358 40432 36414 40488
rect 36634 40568 36690 40624
rect 37646 40604 37648 40624
rect 37648 40604 37700 40624
rect 37700 40604 37702 40624
rect 37646 40568 37702 40604
rect 38198 40468 38200 40488
rect 38200 40468 38252 40488
rect 38252 40468 38254 40488
rect 38198 40432 38254 40468
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 36634 28056 36690 28112
rect 36726 27376 36782 27432
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 40958 38256 41014 38312
rect 38198 24132 38254 24168
rect 38198 24112 38200 24132
rect 38200 24112 38252 24132
rect 38252 24112 38254 24132
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 39762 24148 39764 24168
rect 39764 24148 39816 24168
rect 39816 24148 39818 24168
rect 39762 24112 39818 24148
rect 46754 49000 46810 49056
rect 46846 46960 46902 47016
rect 46846 46280 46902 46336
rect 45742 42200 45798 42256
rect 46846 42880 46902 42936
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 46478 40160 46534 40216
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 45558 23840 45614 23896
rect 46846 33360 46902 33416
rect 46202 26560 46258 26616
rect 45558 17720 45614 17776
rect 46846 29280 46902 29336
rect 46754 21800 46810 21856
rect 47398 38292 47400 38312
rect 47400 38292 47452 38312
rect 47452 38292 47454 38312
rect 47398 38256 47454 38292
rect 48134 44940 48190 44976
rect 48134 44920 48136 44940
rect 48136 44920 48188 44940
rect 48188 44920 48190 44940
rect 48134 41520 48190 41576
rect 48134 39480 48190 39536
rect 48134 38120 48190 38176
rect 48226 37440 48282 37496
rect 48134 36080 48190 36136
rect 48134 32680 48190 32736
rect 48134 28600 48190 28656
rect 48134 27920 48190 27976
rect 48134 25880 48190 25936
rect 48134 22480 48190 22536
rect 48134 20440 48190 20496
rect 48134 19080 48190 19136
rect 48134 17040 48190 17096
rect 48134 15000 48190 15056
rect 48134 13640 48190 13696
rect 48134 12960 48190 13016
rect 46846 12280 46902 12336
rect 47950 8200 48006 8256
rect 46846 2080 46902 2136
rect 48134 6860 48190 6896
rect 48134 6840 48136 6860
rect 48136 6840 48188 6860
rect 48188 6840 48190 6860
rect 48134 5480 48190 5536
rect 48226 1400 48282 1456
rect 46570 40 46626 96
<< metal3 >>
rect 0 49588 800 49828
rect 46749 49058 46815 49061
rect 49200 49058 50000 49148
rect 46749 49056 50000 49058
rect 46749 49000 46754 49056
rect 46810 49000 50000 49056
rect 46749 48998 50000 49000
rect 46749 48995 46815 48998
rect 49200 48908 50000 48998
rect 0 48378 800 48468
rect 3601 48378 3667 48381
rect 0 48376 3667 48378
rect 0 48320 3606 48376
rect 3662 48320 3667 48376
rect 0 48318 3667 48320
rect 0 48228 800 48318
rect 3601 48315 3667 48318
rect 49200 48228 50000 48468
rect 0 47698 800 47788
rect 2773 47698 2839 47701
rect 0 47696 2839 47698
rect 0 47640 2778 47696
rect 2834 47640 2839 47696
rect 0 47638 2839 47640
rect 0 47548 800 47638
rect 2773 47635 2839 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 46841 47018 46907 47021
rect 49200 47018 50000 47108
rect 46841 47016 50000 47018
rect 46841 46960 46846 47016
rect 46902 46960 50000 47016
rect 46841 46958 50000 46960
rect 46841 46955 46907 46958
rect 49200 46868 50000 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 0 46338 800 46428
rect 1669 46338 1735 46341
rect 0 46336 1735 46338
rect 0 46280 1674 46336
rect 1730 46280 1735 46336
rect 0 46278 1735 46280
rect 0 46188 800 46278
rect 1669 46275 1735 46278
rect 46841 46338 46907 46341
rect 49200 46338 50000 46428
rect 46841 46336 50000 46338
rect 46841 46280 46846 46336
rect 46902 46280 50000 46336
rect 46841 46278 50000 46280
rect 46841 46275 46907 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 49200 46188 50000 46278
rect 0 45658 800 45748
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 3693 45658 3759 45661
rect 0 45656 3759 45658
rect 0 45600 3698 45656
rect 3754 45600 3759 45656
rect 0 45598 3759 45600
rect 0 45508 800 45598
rect 3693 45595 3759 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 48129 44978 48195 44981
rect 49200 44978 50000 45068
rect 48129 44976 50000 44978
rect 48129 44920 48134 44976
rect 48190 44920 50000 44976
rect 48129 44918 50000 44920
rect 48129 44915 48195 44918
rect 49200 44828 50000 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 0 44148 800 44388
rect 49200 44148 50000 44388
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 0 43618 800 43708
rect 3969 43618 4035 43621
rect 0 43616 4035 43618
rect 0 43560 3974 43616
rect 4030 43560 4035 43616
rect 0 43558 4035 43560
rect 0 43468 800 43558
rect 3969 43555 4035 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 0 42788 800 43028
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 46841 42938 46907 42941
rect 49200 42938 50000 43028
rect 46841 42936 50000 42938
rect 46841 42880 46846 42936
rect 46902 42880 50000 42936
rect 46841 42878 50000 42880
rect 46841 42875 46907 42878
rect 49200 42788 50000 42878
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 45737 42258 45803 42261
rect 49200 42258 50000 42348
rect 45737 42256 50000 42258
rect 45737 42200 45742 42256
rect 45798 42200 50000 42256
rect 45737 42198 50000 42200
rect 45737 42195 45803 42198
rect 49200 42108 50000 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 0 41578 800 41668
rect 3325 41578 3391 41581
rect 0 41576 3391 41578
rect 0 41520 3330 41576
rect 3386 41520 3391 41576
rect 0 41518 3391 41520
rect 0 41428 800 41518
rect 3325 41515 3391 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41668
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41428 50000 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 33869 41034 33935 41037
rect 34789 41034 34855 41037
rect 33869 41032 34855 41034
rect 0 40898 800 40988
rect 33869 40976 33874 41032
rect 33930 40976 34794 41032
rect 34850 40976 34855 41032
rect 33869 40974 34855 40976
rect 33869 40971 33935 40974
rect 34789 40971 34855 40974
rect 3417 40898 3483 40901
rect 0 40896 3483 40898
rect 0 40840 3422 40896
rect 3478 40840 3483 40896
rect 0 40838 3483 40840
rect 0 40748 800 40838
rect 3417 40835 3483 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 36629 40626 36695 40629
rect 37641 40626 37707 40629
rect 36629 40624 37707 40626
rect 36629 40568 36634 40624
rect 36690 40568 37646 40624
rect 37702 40568 37707 40624
rect 36629 40566 37707 40568
rect 36629 40563 36695 40566
rect 37641 40563 37707 40566
rect 36353 40490 36419 40493
rect 38193 40490 38259 40493
rect 36353 40488 38259 40490
rect 36353 40432 36358 40488
rect 36414 40432 38198 40488
rect 38254 40432 38259 40488
rect 36353 40430 38259 40432
rect 36353 40427 36419 40430
rect 38193 40427 38259 40430
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 46473 40218 46539 40221
rect 49200 40218 50000 40308
rect 46473 40216 50000 40218
rect 46473 40160 46478 40216
rect 46534 40160 50000 40216
rect 46473 40158 50000 40160
rect 46473 40155 46539 40158
rect 49200 40068 50000 40158
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39388 800 39628
rect 48129 39538 48195 39541
rect 49200 39538 50000 39628
rect 48129 39536 50000 39538
rect 48129 39480 48134 39536
rect 48190 39480 50000 39536
rect 48129 39478 50000 39480
rect 48129 39475 48195 39478
rect 49200 39388 50000 39478
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 0 38708 800 38948
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 40953 38314 41019 38317
rect 47393 38314 47459 38317
rect 40953 38312 47459 38314
rect 40953 38256 40958 38312
rect 41014 38256 47398 38312
rect 47454 38256 47459 38312
rect 40953 38254 47459 38256
rect 40953 38251 41019 38254
rect 47393 38251 47459 38254
rect 48129 38178 48195 38181
rect 49200 38178 50000 38268
rect 48129 38176 50000 38178
rect 48129 38120 48134 38176
rect 48190 38120 50000 38176
rect 48129 38118 50000 38120
rect 48129 38115 48195 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 49200 38028 50000 38118
rect 0 37348 800 37588
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 48221 37498 48287 37501
rect 49200 37498 50000 37588
rect 48221 37496 50000 37498
rect 48221 37440 48226 37496
rect 48282 37440 50000 37496
rect 48221 37438 50000 37440
rect 48221 37435 48287 37438
rect 49200 37348 50000 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 0 36668 800 36908
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 35988 800 36228
rect 48129 36138 48195 36141
rect 49200 36138 50000 36228
rect 48129 36136 50000 36138
rect 48129 36080 48134 36136
rect 48190 36080 50000 36136
rect 48129 36078 50000 36080
rect 48129 36075 48195 36078
rect 49200 35988 50000 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 49200 35308 50000 35548
rect 0 34628 800 34868
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 49200 34628 50000 34868
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 33948 800 34188
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 46841 33418 46907 33421
rect 49200 33418 50000 33508
rect 46841 33416 50000 33418
rect 46841 33360 46846 33416
rect 46902 33360 50000 33416
rect 46841 33358 50000 33360
rect 46841 33355 46907 33358
rect 49200 33268 50000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 32305 33146 32371 33149
rect 33133 33146 33199 33149
rect 32305 33144 33199 33146
rect 32305 33088 32310 33144
rect 32366 33088 33138 33144
rect 33194 33088 33199 33144
rect 32305 33086 33199 33088
rect 32305 33083 32371 33086
rect 33133 33083 33199 33086
rect 0 32738 800 32828
rect 2773 32738 2839 32741
rect 0 32736 2839 32738
rect 0 32680 2778 32736
rect 2834 32680 2839 32736
rect 0 32678 2839 32680
rect 0 32588 800 32678
rect 2773 32675 2839 32678
rect 48129 32738 48195 32741
rect 49200 32738 50000 32828
rect 48129 32736 50000 32738
rect 48129 32680 48134 32736
rect 48190 32680 50000 32736
rect 48129 32678 50000 32680
rect 48129 32675 48195 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 49200 32588 50000 32678
rect 0 31908 800 32148
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 49200 31228 50000 31468
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 0 30548 800 30788
rect 49200 30548 50000 30788
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 0 29868 800 30108
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 25589 29610 25655 29613
rect 28073 29610 28139 29613
rect 25589 29608 28139 29610
rect 25589 29552 25594 29608
rect 25650 29552 28078 29608
rect 28134 29552 28139 29608
rect 25589 29550 28139 29552
rect 25589 29547 25655 29550
rect 28073 29547 28139 29550
rect 0 29188 800 29428
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 46841 29338 46907 29341
rect 49200 29338 50000 29428
rect 46841 29336 50000 29338
rect 46841 29280 46846 29336
rect 46902 29280 50000 29336
rect 46841 29278 50000 29280
rect 46841 29275 46907 29278
rect 49200 29188 50000 29278
rect 25773 29066 25839 29069
rect 26141 29066 26207 29069
rect 25773 29064 26207 29066
rect 25773 29008 25778 29064
rect 25834 29008 26146 29064
rect 26202 29008 26207 29064
rect 25773 29006 26207 29008
rect 25773 29003 25839 29006
rect 26141 29003 26207 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 48129 28658 48195 28661
rect 49200 28658 50000 28748
rect 48129 28656 50000 28658
rect 48129 28600 48134 28656
rect 48190 28600 50000 28656
rect 48129 28598 50000 28600
rect 48129 28595 48195 28598
rect 49200 28508 50000 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 31937 28114 32003 28117
rect 36629 28114 36695 28117
rect 31937 28112 36695 28114
rect 0 27828 800 28068
rect 31937 28056 31942 28112
rect 31998 28056 36634 28112
rect 36690 28056 36695 28112
rect 31937 28054 36695 28056
rect 31937 28051 32003 28054
rect 36629 28051 36695 28054
rect 48129 27978 48195 27981
rect 49200 27978 50000 28068
rect 48129 27976 50000 27978
rect 48129 27920 48134 27976
rect 48190 27920 50000 27976
rect 48129 27918 50000 27920
rect 48129 27915 48195 27918
rect 49200 27828 50000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 24117 27434 24183 27437
rect 26509 27434 26575 27437
rect 24117 27432 26575 27434
rect 0 27148 800 27388
rect 24117 27376 24122 27432
rect 24178 27376 26514 27432
rect 26570 27376 26575 27432
rect 24117 27374 26575 27376
rect 24117 27371 24183 27374
rect 26509 27371 26575 27374
rect 30557 27434 30623 27437
rect 36721 27434 36787 27437
rect 30557 27432 36787 27434
rect 30557 27376 30562 27432
rect 30618 27376 36726 27432
rect 36782 27376 36787 27432
rect 30557 27374 36787 27376
rect 30557 27371 30623 27374
rect 36721 27371 36787 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 46197 26618 46263 26621
rect 49200 26618 50000 26708
rect 46197 26616 50000 26618
rect 46197 26560 46202 26616
rect 46258 26560 50000 26616
rect 46197 26558 50000 26560
rect 46197 26555 46263 26558
rect 49200 26468 50000 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 0 25788 800 26028
rect 48129 25938 48195 25941
rect 49200 25938 50000 26028
rect 48129 25936 50000 25938
rect 48129 25880 48134 25936
rect 48190 25880 50000 25936
rect 48129 25878 50000 25880
rect 48129 25875 48195 25878
rect 49200 25788 50000 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25348
rect 2773 25258 2839 25261
rect 0 25256 2839 25258
rect 0 25200 2778 25256
rect 2834 25200 2839 25256
rect 0 25198 2839 25200
rect 0 25108 800 25198
rect 2773 25195 2839 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 49200 24428 50000 24668
rect 38193 24170 38259 24173
rect 39757 24170 39823 24173
rect 38193 24168 39823 24170
rect 38193 24112 38198 24168
rect 38254 24112 39762 24168
rect 39818 24112 39823 24168
rect 38193 24110 39823 24112
rect 38193 24107 38259 24110
rect 39757 24107 39823 24110
rect 0 23898 800 23988
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 2773 23898 2839 23901
rect 0 23896 2839 23898
rect 0 23840 2778 23896
rect 2834 23840 2839 23896
rect 0 23838 2839 23840
rect 0 23748 800 23838
rect 2773 23835 2839 23838
rect 45553 23898 45619 23901
rect 49200 23898 50000 23988
rect 45553 23896 50000 23898
rect 45553 23840 45558 23896
rect 45614 23840 50000 23896
rect 45553 23838 50000 23840
rect 45553 23835 45619 23838
rect 49200 23748 50000 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23068 800 23308
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 48129 22538 48195 22541
rect 49200 22538 50000 22628
rect 48129 22536 50000 22538
rect 48129 22480 48134 22536
rect 48190 22480 50000 22536
rect 48129 22478 50000 22480
rect 48129 22475 48195 22478
rect 49200 22388 50000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 0 21858 800 21948
rect 2773 21858 2839 21861
rect 0 21856 2839 21858
rect 0 21800 2778 21856
rect 2834 21800 2839 21856
rect 0 21798 2839 21800
rect 0 21708 800 21798
rect 2773 21795 2839 21798
rect 46749 21858 46815 21861
rect 49200 21858 50000 21948
rect 46749 21856 50000 21858
rect 46749 21800 46754 21856
rect 46810 21800 50000 21856
rect 46749 21798 50000 21800
rect 46749 21795 46815 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 49200 21708 50000 21798
rect 0 21028 800 21268
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 0 20498 800 20588
rect 2773 20498 2839 20501
rect 0 20496 2839 20498
rect 0 20440 2778 20496
rect 2834 20440 2839 20496
rect 0 20438 2839 20440
rect 0 20348 800 20438
rect 2773 20435 2839 20438
rect 48129 20498 48195 20501
rect 49200 20498 50000 20588
rect 48129 20496 50000 20498
rect 48129 20440 48134 20496
rect 48190 20440 50000 20496
rect 48129 20438 50000 20440
rect 48129 20435 48195 20438
rect 49200 20348 50000 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 49200 19668 50000 19908
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 0 18988 800 19228
rect 48129 19138 48195 19141
rect 49200 19138 50000 19228
rect 48129 19136 50000 19138
rect 48129 19080 48134 19136
rect 48190 19080 50000 19136
rect 48129 19078 50000 19080
rect 48129 19075 48195 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 49200 18988 50000 19078
rect 0 18458 800 18548
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 2773 18458 2839 18461
rect 0 18456 2839 18458
rect 0 18400 2778 18456
rect 2834 18400 2839 18456
rect 0 18398 2839 18400
rect 0 18308 800 18398
rect 2773 18395 2839 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 45553 17778 45619 17781
rect 49200 17778 50000 17868
rect 45553 17776 50000 17778
rect 45553 17720 45558 17776
rect 45614 17720 50000 17776
rect 45553 17718 50000 17720
rect 45553 17715 45619 17718
rect 49200 17628 50000 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 0 17098 800 17188
rect 2773 17098 2839 17101
rect 0 17096 2839 17098
rect 0 17040 2778 17096
rect 2834 17040 2839 17096
rect 0 17038 2839 17040
rect 0 16948 800 17038
rect 2773 17035 2839 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17188
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 16948 50000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 0 16268 800 16508
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 49200 15588 50000 15828
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 0 15058 800 15148
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14908 800 14998
rect 2773 14995 2839 14998
rect 48129 15058 48195 15061
rect 49200 15058 50000 15148
rect 48129 15056 50000 15058
rect 48129 15000 48134 15056
rect 48190 15000 50000 15056
rect 48129 14998 50000 15000
rect 48129 14995 48195 14998
rect 49200 14908 50000 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 0 14378 800 14468
rect 2773 14378 2839 14381
rect 0 14376 2839 14378
rect 0 14320 2778 14376
rect 2834 14320 2839 14376
rect 0 14318 2839 14320
rect 0 14228 800 14318
rect 2773 14315 2839 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 0 13548 800 13788
rect 48129 13698 48195 13701
rect 49200 13698 50000 13788
rect 48129 13696 50000 13698
rect 48129 13640 48134 13696
rect 48190 13640 50000 13696
rect 48129 13638 50000 13640
rect 48129 13635 48195 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 49200 13548 50000 13638
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 48129 13018 48195 13021
rect 49200 13018 50000 13108
rect 48129 13016 50000 13018
rect 48129 12960 48134 13016
rect 48190 12960 50000 13016
rect 48129 12958 50000 12960
rect 48129 12955 48195 12958
rect 49200 12868 50000 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12188 800 12428
rect 46841 12338 46907 12341
rect 49200 12338 50000 12428
rect 46841 12336 50000 12338
rect 46841 12280 46846 12336
rect 46902 12280 50000 12336
rect 46841 12278 50000 12280
rect 46841 12275 46907 12278
rect 49200 12188 50000 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 0 11658 800 11748
rect 2773 11658 2839 11661
rect 0 11656 2839 11658
rect 0 11600 2778 11656
rect 2834 11600 2839 11656
rect 0 11598 2839 11600
rect 0 11508 800 11598
rect 2773 11595 2839 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 49200 10828 50000 11068
rect 0 10298 800 10388
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 3233 10298 3299 10301
rect 0 10296 3299 10298
rect 0 10240 3238 10296
rect 3294 10240 3299 10296
rect 0 10238 3299 10240
rect 0 10148 800 10238
rect 3233 10235 3299 10238
rect 49200 10148 50000 10388
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 0 9618 800 9708
rect 2865 9618 2931 9621
rect 0 9616 2931 9618
rect 0 9560 2870 9616
rect 2926 9560 2931 9616
rect 0 9558 2931 9560
rect 0 9468 800 9558
rect 2865 9555 2931 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 49200 8788 50000 9028
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 0 8108 800 8348
rect 47945 8258 48011 8261
rect 49200 8258 50000 8348
rect 47945 8256 50000 8258
rect 47945 8200 47950 8256
rect 48006 8200 50000 8256
rect 47945 8198 50000 8200
rect 47945 8195 48011 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 49200 8108 50000 8198
rect 0 7578 800 7668
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 2773 7578 2839 7581
rect 0 7576 2839 7578
rect 0 7520 2778 7576
rect 2834 7520 2839 7576
rect 0 7518 2839 7520
rect 0 7428 800 7518
rect 2773 7515 2839 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6988
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6748 800 6838
rect 2773 6835 2839 6838
rect 48129 6898 48195 6901
rect 49200 6898 50000 6988
rect 48129 6896 50000 6898
rect 48129 6840 48134 6896
rect 48190 6840 50000 6896
rect 48129 6838 50000 6840
rect 48129 6835 48195 6838
rect 49200 6748 50000 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 49200 6068 50000 6308
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 0 5538 800 5628
rect 2865 5538 2931 5541
rect 0 5536 2931 5538
rect 0 5480 2870 5536
rect 2926 5480 2931 5536
rect 0 5478 2931 5480
rect 0 5388 800 5478
rect 2865 5475 2931 5478
rect 48129 5538 48195 5541
rect 49200 5538 50000 5628
rect 48129 5536 50000 5538
rect 48129 5480 48134 5536
rect 48190 5480 50000 5536
rect 48129 5478 50000 5480
rect 48129 5475 48195 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 49200 5388 50000 5478
rect 0 4858 800 4948
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 3141 4858 3207 4861
rect 0 4856 3207 4858
rect 0 4800 3146 4856
rect 3202 4800 3207 4856
rect 0 4798 3207 4800
rect 0 4708 800 4798
rect 3141 4795 3207 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 49200 4028 50000 4268
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 0 3498 800 3588
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3348 800 3438
rect 1853 3435 1919 3438
rect 49200 3348 50000 3588
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 0 2818 800 2908
rect 4061 2818 4127 2821
rect 0 2816 4127 2818
rect 0 2760 4066 2816
rect 4122 2760 4127 2816
rect 0 2758 4127 2760
rect 0 2668 800 2758
rect 4061 2755 4127 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 46841 2138 46907 2141
rect 49200 2138 50000 2228
rect 46841 2136 50000 2138
rect 46841 2080 46846 2136
rect 46902 2080 50000 2136
rect 46841 2078 50000 2080
rect 46841 2075 46907 2078
rect 49200 1988 50000 2078
rect 0 1458 800 1548
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1308 800 1398
rect 2773 1395 2839 1398
rect 48221 1458 48287 1461
rect 49200 1458 50000 1548
rect 48221 1456 50000 1458
rect 48221 1400 48226 1456
rect 48282 1400 50000 1456
rect 48221 1398 50000 1400
rect 48221 1395 48287 1398
rect 49200 1308 50000 1398
rect 0 628 800 868
rect 46565 98 46631 101
rect 49200 98 50000 188
rect 46565 96 50000 98
rect 46565 40 46570 96
rect 46626 40 50000 96
rect 46565 38 50000 40
rect 46565 35 46631 38
rect 49200 -52 50000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22724 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1649977179
transform 1 0 27600 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1649977179
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106
timestamp 1649977179
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_205
timestamp 1649977179
transform 1 0 19964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1649977179
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_263
timestamp 1649977179
transform 1 0 25300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1649977179
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1649977179
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1649977179
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1649977179
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1649977179
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1649977179
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1649977179
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1649977179
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1649977179
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_470
timestamp 1649977179
transform 1 0 44344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1649977179
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_508 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_94
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1649977179
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_121
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_126
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_155
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_260
timestamp 1649977179
transform 1 0 25024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_267
timestamp 1649977179
transform 1 0 25668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_302
timestamp 1649977179
transform 1 0 28888 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_314
timestamp 1649977179
transform 1 0 29992 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_326
timestamp 1649977179
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1649977179
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_358
timestamp 1649977179
transform 1 0 34040 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_370
timestamp 1649977179
transform 1 0 35144 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1649977179
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1649977179
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_428
timestamp 1649977179
transform 1 0 40480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_435
timestamp 1649977179
transform 1 0 41124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1649977179
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_470
timestamp 1649977179
transform 1 0 44344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1649977179
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1649977179
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_95
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_144
timestamp 1649977179
transform 1 0 14352 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_156
timestamp 1649977179
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_168
timestamp 1649977179
transform 1 0 16560 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_174
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_230
timestamp 1649977179
transform 1 0 22264 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_242
timestamp 1649977179
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1649977179
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_261
timestamp 1649977179
transform 1 0 25116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_284
timestamp 1649977179
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_291
timestamp 1649977179
transform 1 0 27876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_298
timestamp 1649977179
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1649977179
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_329
timestamp 1649977179
transform 1 0 31372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_334
timestamp 1649977179
transform 1 0 31832 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_341
timestamp 1649977179
transform 1 0 32476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_353
timestamp 1649977179
transform 1 0 33580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp 1649977179
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1649977179
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_442
timestamp 1649977179
transform 1 0 41768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_467
timestamp 1649977179
transform 1 0 44068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1649977179
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1649977179
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1649977179
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp 1649977179
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_40
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_48
timestamp 1649977179
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1649977179
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_64
timestamp 1649977179
transform 1 0 6992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_68
timestamp 1649977179
transform 1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_101
timestamp 1649977179
transform 1 0 10396 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1649977179
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_155
timestamp 1649977179
transform 1 0 15364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1649977179
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_212
timestamp 1649977179
transform 1 0 20608 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_231
timestamp 1649977179
transform 1 0 22356 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_243
timestamp 1649977179
transform 1 0 23460 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_255
timestamp 1649977179
transform 1 0 24564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_263
timestamp 1649977179
transform 1 0 25300 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_267
timestamp 1649977179
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_411
timestamp 1649977179
transform 1 0 38916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_418
timestamp 1649977179
transform 1 0 39560 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_422
timestamp 1649977179
transform 1 0 39928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_426
timestamp 1649977179
transform 1 0 40296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_430
timestamp 1649977179
transform 1 0 40664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_434
timestamp 1649977179
transform 1 0 41032 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_440
timestamp 1649977179
transform 1 0 41584 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1649977179
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_452
timestamp 1649977179
transform 1 0 42688 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_460
timestamp 1649977179
transform 1 0 43424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_464
timestamp 1649977179
transform 1 0 43792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_471
timestamp 1649977179
transform 1 0 44436 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1649977179
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_508
timestamp 1649977179
transform 1 0 47840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1649977179
transform 1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 1649977179
transform 1 0 2576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_33
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1649977179
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_44
timestamp 1649977179
transform 1 0 5152 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_52
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_58
timestamp 1649977179
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_70
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1649977179
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_88
timestamp 1649977179
transform 1 0 9200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_100
timestamp 1649977179
transform 1 0 10304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_112
timestamp 1649977179
transform 1 0 11408 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_124
timestamp 1649977179
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_200
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_207
timestamp 1649977179
transform 1 0 20148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_219
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_231
timestamp 1649977179
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1649977179
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_449
timestamp 1649977179
transform 1 0 42412 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_461
timestamp 1649977179
transform 1 0 43516 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_472
timestamp 1649977179
transform 1 0 44528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_483
timestamp 1649977179
transform 1 0 45540 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1649977179
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_10
timestamp 1649977179
transform 1 0 2024 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_469
timestamp 1649977179
transform 1 0 44252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_475
timestamp 1649977179
transform 1 0 44804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1649977179
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_508
timestamp 1649977179
transform 1 0 47840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 1649977179
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_17
timestamp 1649977179
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1649977179
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_44
timestamp 1649977179
transform 1 0 5152 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_56
timestamp 1649977179
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_68
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_483
timestamp 1649977179
transform 1 0 45540 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_487
timestamp 1649977179
transform 1 0 45908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1649977179
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_32
timestamp 1649977179
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1649977179
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_489
timestamp 1649977179
transform 1 0 46092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_493
timestamp 1649977179
transform 1 0 46460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_500
timestamp 1649977179
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_508
timestamp 1649977179
transform 1 0 47840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_11
timestamp 1649977179
transform 1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_17
timestamp 1649977179
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1649977179
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1649977179
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1649977179
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1649977179
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1649977179
transform 1 0 47840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1649977179
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1649977179
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_32
timestamp 1649977179
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1649977179
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_14
timestamp 1649977179
transform 1 0 2392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_14
timestamp 1649977179
transform 1 0 2392 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1649977179
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1649977179
transform 1 0 2392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1649977179
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_32
timestamp 1649977179
transform 1 0 4048 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_44
timestamp 1649977179
transform 1 0 5152 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_56
timestamp 1649977179
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_68
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_207
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_219
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_231
timestamp 1649977179
transform 1 0 22356 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_243
timestamp 1649977179
transform 1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_273
timestamp 1649977179
transform 1 0 26220 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_278
timestamp 1649977179
transform 1 0 26680 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_290
timestamp 1649977179
transform 1 0 27784 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_302
timestamp 1649977179
transform 1 0 28888 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_32
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1649977179
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1649977179
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_16
timestamp 1649977179
transform 1 0 2576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1649977179
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1649977179
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_31
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1649977179
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_493
timestamp 1649977179
transform 1 0 46460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_499
timestamp 1649977179
transform 1 0 47012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1649977179
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_14
timestamp 1649977179
transform 1 0 2392 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_512
timestamp 1649977179
transform 1 0 48208 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_489
timestamp 1649977179
transform 1 0 46092 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_493
timestamp 1649977179
transform 1 0 46460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_500
timestamp 1649977179
transform 1 0 47104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_508
timestamp 1649977179
transform 1 0 47840 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_512
timestamp 1649977179
transform 1 0 48208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_32
timestamp 1649977179
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1649977179
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_508
timestamp 1649977179
transform 1 0 47840 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_32
timestamp 1649977179
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_44
timestamp 1649977179
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_68
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_512
timestamp 1649977179
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_32
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_44
timestamp 1649977179
transform 1 0 5152 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_508
timestamp 1649977179
transform 1 0 47840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_14
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_507
timestamp 1649977179
transform 1 0 47748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_515
timestamp 1649977179
transform 1 0 48484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_513
timestamp 1649977179
transform 1 0 48300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_11
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_17
timestamp 1649977179
transform 1 0 2668 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1649977179
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_427
timestamp 1649977179
transform 1 0 40388 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_439
timestamp 1649977179
transform 1 0 41492 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_451
timestamp 1649977179
transform 1 0 42596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_463
timestamp 1649977179
transform 1 0 43700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1649977179
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_32
timestamp 1649977179
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_44
timestamp 1649977179
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_421
timestamp 1649977179
transform 1 0 39836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_436
timestamp 1649977179
transform 1 0 41216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_456
timestamp 1649977179
transform 1 0 43056 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_464
timestamp 1649977179
transform 1 0 43792 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_470
timestamp 1649977179
transform 1 0 44344 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_482
timestamp 1649977179
transform 1 0 45448 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_494
timestamp 1649977179
transform 1 0 46552 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1649977179
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1649977179
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_14
timestamp 1649977179
transform 1 0 2392 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_129
timestamp 1649977179
transform 1 0 12972 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_404
timestamp 1649977179
transform 1 0 38272 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_415
timestamp 1649977179
transform 1 0 39284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_430
timestamp 1649977179
transform 1 0 40664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_439
timestamp 1649977179
transform 1 0 41492 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_447
timestamp 1649977179
transform 1 0 42228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_468
timestamp 1649977179
transform 1 0 44160 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1649977179
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1649977179
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_130
timestamp 1649977179
transform 1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_155
timestamp 1649977179
transform 1 0 15364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_453
timestamp 1649977179
transform 1 0 42780 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_465
timestamp 1649977179
transform 1 0 43884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_469
timestamp 1649977179
transform 1 0 44252 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_478
timestamp 1649977179
transform 1 0 45080 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_489
timestamp 1649977179
transform 1 0 46092 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1649977179
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_508
timestamp 1649977179
transform 1 0 47840 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_14
timestamp 1649977179
transform 1 0 2392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1649977179
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_411
timestamp 1649977179
transform 1 0 38916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_430
timestamp 1649977179
transform 1 0 40664 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_448
timestamp 1649977179
transform 1 0 42320 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_456
timestamp 1649977179
transform 1 0 43056 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_463
timestamp 1649977179
transform 1 0 43700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1649977179
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_487
timestamp 1649977179
transform 1 0 45908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1649977179
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_285
timestamp 1649977179
transform 1 0 27324 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_297
timestamp 1649977179
transform 1 0 28428 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_309
timestamp 1649977179
transform 1 0 29532 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_321
timestamp 1649977179
transform 1 0 30636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1649977179
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_342
timestamp 1649977179
transform 1 0 32568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_346
timestamp 1649977179
transform 1 0 32936 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_363
timestamp 1649977179
transform 1 0 34500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_375
timestamp 1649977179
transform 1 0 35604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1649977179
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_409
timestamp 1649977179
transform 1 0 38732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_416
timestamp 1649977179
transform 1 0 39376 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_424
timestamp 1649977179
transform 1 0 40112 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_433
timestamp 1649977179
transform 1 0 40940 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_439
timestamp 1649977179
transform 1 0 41492 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_444
timestamp 1649977179
transform 1 0 41952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_452
timestamp 1649977179
transform 1 0 42688 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_468
timestamp 1649977179
transform 1 0 44160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_480
timestamp 1649977179
transform 1 0 45264 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_500
timestamp 1649977179
transform 1 0 47104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1649977179
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 1649977179
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_257
timestamp 1649977179
transform 1 0 24748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_274
timestamp 1649977179
transform 1 0 26312 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_294
timestamp 1649977179
transform 1 0 28152 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1649977179
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_315
timestamp 1649977179
transform 1 0 30084 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_320
timestamp 1649977179
transform 1 0 30544 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_332
timestamp 1649977179
transform 1 0 31648 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_349
timestamp 1649977179
transform 1 0 33212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_370
timestamp 1649977179
transform 1 0 35144 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_378
timestamp 1649977179
transform 1 0 35880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_396
timestamp 1649977179
transform 1 0 37536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_404
timestamp 1649977179
transform 1 0 38272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_408
timestamp 1649977179
transform 1 0 38640 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_412
timestamp 1649977179
transform 1 0 39008 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_441
timestamp 1649977179
transform 1 0 41676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_461
timestamp 1649977179
transform 1 0 43516 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_467
timestamp 1649977179
transform 1 0 44068 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1649977179
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_485
timestamp 1649977179
transform 1 0 45724 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1649977179
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1649977179
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1649977179
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1649977179
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_290
timestamp 1649977179
transform 1 0 27784 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_298
timestamp 1649977179
transform 1 0 28520 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_310
timestamp 1649977179
transform 1 0 29624 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_345
timestamp 1649977179
transform 1 0 32844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_351
timestamp 1649977179
transform 1 0 33396 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_371
timestamp 1649977179
transform 1 0 35236 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_378
timestamp 1649977179
transform 1 0 35880 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1649977179
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_401
timestamp 1649977179
transform 1 0 37996 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_409
timestamp 1649977179
transform 1 0 38732 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_479
timestamp 1649977179
transform 1 0 45172 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_491
timestamp 1649977179
transform 1 0 46276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_508
timestamp 1649977179
transform 1 0 47840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_11
timestamp 1649977179
transform 1 0 2116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_16
timestamp 1649977179
transform 1 0 2576 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1649977179
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_269
timestamp 1649977179
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_276
timestamp 1649977179
transform 1 0 26496 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_284
timestamp 1649977179
transform 1 0 27232 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1649977179
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1649977179
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_336
timestamp 1649977179
transform 1 0 32016 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_348
timestamp 1649977179
transform 1 0 33120 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_358
timestamp 1649977179
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_371
timestamp 1649977179
transform 1 0 35236 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_378
timestamp 1649977179
transform 1 0 35880 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_390
timestamp 1649977179
transform 1 0 36984 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_394
timestamp 1649977179
transform 1 0 37352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_403
timestamp 1649977179
transform 1 0 38180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_411
timestamp 1649977179
transform 1 0 38916 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_416
timestamp 1649977179
transform 1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_428
timestamp 1649977179
transform 1 0 40480 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_440
timestamp 1649977179
transform 1 0 41584 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_452
timestamp 1649977179
transform 1 0 42688 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_458
timestamp 1649977179
transform 1 0 43240 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_470
timestamp 1649977179
transform 1 0 44344 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_480
timestamp 1649977179
transform 1 0 45264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_492
timestamp 1649977179
transform 1 0 46368 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1649977179
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_9
timestamp 1649977179
transform 1 0 1932 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1649977179
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1649977179
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1649977179
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_263
timestamp 1649977179
transform 1 0 25300 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1649977179
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_286
timestamp 1649977179
transform 1 0 27416 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1649977179
transform 1 0 28244 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_302
timestamp 1649977179
transform 1 0 28888 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_314
timestamp 1649977179
transform 1 0 29992 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_321
timestamp 1649977179
transform 1 0 30636 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_365
timestamp 1649977179
transform 1 0 34684 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_377
timestamp 1649977179
transform 1 0 35788 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_384
timestamp 1649977179
transform 1 0 36432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_401
timestamp 1649977179
transform 1 0 37996 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_413
timestamp 1649977179
transform 1 0 39100 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_426
timestamp 1649977179
transform 1 0 40296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_438
timestamp 1649977179
transform 1 0 41400 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_444
timestamp 1649977179
transform 1 0 41952 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_457
timestamp 1649977179
transform 1 0 43148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_465
timestamp 1649977179
transform 1 0 43884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_489
timestamp 1649977179
transform 1 0 46092 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1649977179
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1649977179
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_14
timestamp 1649977179
transform 1 0 2392 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1649977179
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_269
timestamp 1649977179
transform 1 0 25852 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_278
timestamp 1649977179
transform 1 0 26680 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_286
timestamp 1649977179
transform 1 0 27416 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_298
timestamp 1649977179
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1649977179
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_313
timestamp 1649977179
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_320
timestamp 1649977179
transform 1 0 30544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1649977179
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_335
timestamp 1649977179
transform 1 0 31924 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_349
timestamp 1649977179
transform 1 0 33212 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1649977179
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_393
timestamp 1649977179
transform 1 0 37260 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_405
timestamp 1649977179
transform 1 0 38364 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1649977179
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_430
timestamp 1649977179
transform 1 0 40664 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_438
timestamp 1649977179
transform 1 0 41400 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_450
timestamp 1649977179
transform 1 0 42504 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_484
timestamp 1649977179
transform 1 0 45632 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_490
timestamp 1649977179
transform 1 0 46184 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1649977179
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_257
timestamp 1649977179
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1649977179
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1649977179
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_325
timestamp 1649977179
transform 1 0 31004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1649977179
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_343
timestamp 1649977179
transform 1 0 32660 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_363
timestamp 1649977179
transform 1 0 34500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_375
timestamp 1649977179
transform 1 0 35604 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_382
timestamp 1649977179
transform 1 0 36248 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1649977179
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_396
timestamp 1649977179
transform 1 0 37536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1649977179
transform 1 0 38180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_407
timestamp 1649977179
transform 1 0 38548 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_411
timestamp 1649977179
transform 1 0 38916 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_422
timestamp 1649977179
transform 1 0 39928 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_435
timestamp 1649977179
transform 1 0 41124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_465
timestamp 1649977179
transform 1 0 43884 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_477
timestamp 1649977179
transform 1 0 44988 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1649977179
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_508
timestamp 1649977179
transform 1 0 47840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_11
timestamp 1649977179
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_16
timestamp 1649977179
transform 1 0 2576 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_260
timestamp 1649977179
transform 1 0 25024 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_272
timestamp 1649977179
transform 1 0 26128 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_291
timestamp 1649977179
transform 1 0 27876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_295
timestamp 1649977179
transform 1 0 28244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1649977179
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_317
timestamp 1649977179
transform 1 0 30268 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_323
timestamp 1649977179
transform 1 0 30820 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_347
timestamp 1649977179
transform 1 0 33028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1649977179
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_375
timestamp 1649977179
transform 1 0 35604 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_385
timestamp 1649977179
transform 1 0 36524 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_397
timestamp 1649977179
transform 1 0 37628 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_424
timestamp 1649977179
transform 1 0 40112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_428
timestamp 1649977179
transform 1 0 40480 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_438
timestamp 1649977179
transform 1 0 41400 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_450
timestamp 1649977179
transform 1 0 42504 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_462
timestamp 1649977179
transform 1 0 43608 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1649977179
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_480
timestamp 1649977179
transform 1 0 45264 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_492
timestamp 1649977179
transform 1 0 46368 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_511
timestamp 1649977179
transform 1 0 48116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_515
timestamp 1649977179
transform 1 0 48484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_9
timestamp 1649977179
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_31
timestamp 1649977179
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_43
timestamp 1649977179
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_245
timestamp 1649977179
transform 1 0 23644 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_260
timestamp 1649977179
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1649977179
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_290
timestamp 1649977179
transform 1 0 27784 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_298
timestamp 1649977179
transform 1 0 28520 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_319
timestamp 1649977179
transform 1 0 30452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1649977179
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_357
timestamp 1649977179
transform 1 0 33948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_377
timestamp 1649977179
transform 1 0 35788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_386
timestamp 1649977179
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_411
timestamp 1649977179
transform 1 0 38916 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_419
timestamp 1649977179
transform 1 0 39652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_427
timestamp 1649977179
transform 1 0 40388 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_444
timestamp 1649977179
transform 1 0 41952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_455
timestamp 1649977179
transform 1 0 42964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_459
timestamp 1649977179
transform 1 0 43332 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_470
timestamp 1649977179
transform 1 0 44344 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_482
timestamp 1649977179
transform 1 0 45448 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_492
timestamp 1649977179
transform 1 0 46368 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_496
timestamp 1649977179
transform 1 0 46736 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1649977179
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_508
timestamp 1649977179
transform 1 0 47840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_14
timestamp 1649977179
transform 1 0 2392 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1649977179
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_230
timestamp 1649977179
transform 1 0 22264 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_236
timestamp 1649977179
transform 1 0 22816 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 1649977179
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_269
timestamp 1649977179
transform 1 0 25852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_281
timestamp 1649977179
transform 1 0 26956 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_287
timestamp 1649977179
transform 1 0 27508 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_293
timestamp 1649977179
transform 1 0 28060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1649977179
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_317
timestamp 1649977179
transform 1 0 30268 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_327
timestamp 1649977179
transform 1 0 31188 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_335
timestamp 1649977179
transform 1 0 31924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_343
timestamp 1649977179
transform 1 0 32660 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_350
timestamp 1649977179
transform 1 0 33304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_358
timestamp 1649977179
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_370
timestamp 1649977179
transform 1 0 35144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_390
timestamp 1649977179
transform 1 0 36984 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_398
timestamp 1649977179
transform 1 0 37720 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_404
timestamp 1649977179
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_424
timestamp 1649977179
transform 1 0 40112 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_463
timestamp 1649977179
transform 1 0 43700 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_467
timestamp 1649977179
transform 1 0 44068 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_483
timestamp 1649977179
transform 1 0 45540 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1649977179
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_32
timestamp 1649977179
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1649977179
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_79
timestamp 1649977179
transform 1 0 8372 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_91
timestamp 1649977179
transform 1 0 9476 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_103
timestamp 1649977179
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_248
timestamp 1649977179
transform 1 0 23920 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_256
timestamp 1649977179
transform 1 0 24656 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_260
timestamp 1649977179
transform 1 0 25024 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_272
timestamp 1649977179
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_287
timestamp 1649977179
transform 1 0 27508 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_295
timestamp 1649977179
transform 1 0 28244 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_302
timestamp 1649977179
transform 1 0 28888 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_314
timestamp 1649977179
transform 1 0 29992 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_322
timestamp 1649977179
transform 1 0 30728 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1649977179
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_360
timestamp 1649977179
transform 1 0 34224 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_372
timestamp 1649977179
transform 1 0 35328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_380
timestamp 1649977179
transform 1 0 36064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1649977179
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_424
timestamp 1649977179
transform 1 0 40112 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_436
timestamp 1649977179
transform 1 0 41216 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_465
timestamp 1649977179
transform 1 0 43884 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_475
timestamp 1649977179
transform 1 0 44804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_486
timestamp 1649977179
transform 1 0 45816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_494
timestamp 1649977179
transform 1 0 46552 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_502
timestamp 1649977179
transform 1 0 47288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1649977179
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_12
timestamp 1649977179
transform 1 0 2208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1649977179
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1649977179
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_228
timestamp 1649977179
transform 1 0 22080 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_237
timestamp 1649977179
transform 1 0 22908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1649977179
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_267
timestamp 1649977179
transform 1 0 25668 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_274
timestamp 1649977179
transform 1 0 26312 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_286
timestamp 1649977179
transform 1 0 27416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_290
timestamp 1649977179
transform 1 0 27784 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_294
timestamp 1649977179
transform 1 0 28152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1649977179
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_312
timestamp 1649977179
transform 1 0 29808 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_320
timestamp 1649977179
transform 1 0 30544 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_338
timestamp 1649977179
transform 1 0 32200 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_350
timestamp 1649977179
transform 1 0 33304 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1649977179
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_380
timestamp 1649977179
transform 1 0 36064 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_392
timestamp 1649977179
transform 1 0 37168 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_404
timestamp 1649977179
transform 1 0 38272 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1649977179
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_429
timestamp 1649977179
transform 1 0 40572 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_436
timestamp 1649977179
transform 1 0 41216 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_448
timestamp 1649977179
transform 1 0 42320 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_460
timestamp 1649977179
transform 1 0 43424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_464
timestamp 1649977179
transform 1 0 43792 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_472
timestamp 1649977179
transform 1 0 44528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_483
timestamp 1649977179
transform 1 0 45540 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1649977179
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_73
timestamp 1649977179
transform 1 0 7820 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_83
timestamp 1649977179
transform 1 0 8740 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_96
timestamp 1649977179
transform 1 0 9936 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1649977179
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_234
timestamp 1649977179
transform 1 0 22632 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_246
timestamp 1649977179
transform 1 0 23736 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1649977179
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_284
timestamp 1649977179
transform 1 0 27232 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1649977179
transform 1 0 28244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_314
timestamp 1649977179
transform 1 0 29992 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_347
timestamp 1649977179
transform 1 0 33028 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_356
timestamp 1649977179
transform 1 0 33856 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_368
timestamp 1649977179
transform 1 0 34960 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_380
timestamp 1649977179
transform 1 0 36064 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_387
timestamp 1649977179
transform 1 0 36708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_411
timestamp 1649977179
transform 1 0 38916 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_432
timestamp 1649977179
transform 1 0 40848 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_444
timestamp 1649977179
transform 1 0 41952 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_468
timestamp 1649977179
transform 1 0 44160 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_478
timestamp 1649977179
transform 1 0 45080 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_487
timestamp 1649977179
transform 1 0 45908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_494
timestamp 1649977179
transform 1 0 46552 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_502
timestamp 1649977179
transform 1 0 47288 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_508
timestamp 1649977179
transform 1 0 47840 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1649977179
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_175
timestamp 1649977179
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1649977179
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_241
timestamp 1649977179
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1649977179
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_272
timestamp 1649977179
transform 1 0 26128 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_281
timestamp 1649977179
transform 1 0 26956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_293
timestamp 1649977179
transform 1 0 28060 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_302
timestamp 1649977179
transform 1 0 28888 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_355
timestamp 1649977179
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_370
timestamp 1649977179
transform 1 0 35144 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_380
timestamp 1649977179
transform 1 0 36064 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_400
timestamp 1649977179
transform 1 0 37904 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_408
timestamp 1649977179
transform 1 0 38640 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_439
timestamp 1649977179
transform 1 0 41492 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_460
timestamp 1649977179
transform 1 0 43424 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_472
timestamp 1649977179
transform 1 0 44528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_485
timestamp 1649977179
transform 1 0 45724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_510
timestamp 1649977179
transform 1 0 48024 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_76
timestamp 1649977179
transform 1 0 8096 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_88
timestamp 1649977179
transform 1 0 9200 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_100
timestamp 1649977179
transform 1 0 10304 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_180
timestamp 1649977179
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_190
timestamp 1649977179
transform 1 0 18584 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_202
timestamp 1649977179
transform 1 0 19688 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1649977179
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1649977179
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_245
timestamp 1649977179
transform 1 0 23644 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_253
timestamp 1649977179
transform 1 0 24380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_262
timestamp 1649977179
transform 1 0 25208 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_268
timestamp 1649977179
transform 1 0 25760 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1649977179
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_289
timestamp 1649977179
transform 1 0 27692 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_295
timestamp 1649977179
transform 1 0 28244 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_303
timestamp 1649977179
transform 1 0 28980 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_315
timestamp 1649977179
transform 1 0 30084 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_327
timestamp 1649977179
transform 1 0 31188 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_357
timestamp 1649977179
transform 1 0 33948 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_375
timestamp 1649977179
transform 1 0 35604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1649977179
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_397
timestamp 1649977179
transform 1 0 37628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_437
timestamp 1649977179
transform 1 0 41308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_445
timestamp 1649977179
transform 1 0 42044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_456
timestamp 1649977179
transform 1 0 43056 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_480
timestamp 1649977179
transform 1 0 45264 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_486
timestamp 1649977179
transform 1 0 45816 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_490
timestamp 1649977179
transform 1 0 46184 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_496
timestamp 1649977179
transform 1 0 46736 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_500
timestamp 1649977179
transform 1 0 47104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_508
timestamp 1649977179
transform 1 0 47840 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_159
timestamp 1649977179
transform 1 0 15732 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_164
timestamp 1649977179
transform 1 0 16192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_179
timestamp 1649977179
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1649977179
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_266
timestamp 1649977179
transform 1 0 25576 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_270
timestamp 1649977179
transform 1 0 25944 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_274
timestamp 1649977179
transform 1 0 26312 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_286
timestamp 1649977179
transform 1 0 27416 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_298
timestamp 1649977179
transform 1 0 28520 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1649977179
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_314
timestamp 1649977179
transform 1 0 29992 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_322
timestamp 1649977179
transform 1 0 30728 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_339
timestamp 1649977179
transform 1 0 32292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_351
timestamp 1649977179
transform 1 0 33396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_355
timestamp 1649977179
transform 1 0 33764 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_359
timestamp 1649977179
transform 1 0 34132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_369
timestamp 1649977179
transform 1 0 35052 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_376
timestamp 1649977179
transform 1 0 35696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_388
timestamp 1649977179
transform 1 0 36800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_396
timestamp 1649977179
transform 1 0 37536 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_407
timestamp 1649977179
transform 1 0 38548 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_415
timestamp 1649977179
transform 1 0 39284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_425
timestamp 1649977179
transform 1 0 40204 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_434
timestamp 1649977179
transform 1 0 41032 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_454
timestamp 1649977179
transform 1 0 42872 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_462
timestamp 1649977179
transform 1 0 43608 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_474
timestamp 1649977179
transform 1 0 44712 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_512
timestamp 1649977179
transform 1 0 48208 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_176
timestamp 1649977179
transform 1 0 17296 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_189
timestamp 1649977179
transform 1 0 18492 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_201
timestamp 1649977179
transform 1 0 19596 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1649977179
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1649977179
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_229
timestamp 1649977179
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_247
timestamp 1649977179
transform 1 0 23828 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1649977179
transform 1 0 24932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_265
timestamp 1649977179
transform 1 0 25484 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1649977179
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_286
timestamp 1649977179
transform 1 0 27416 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_294
timestamp 1649977179
transform 1 0 28152 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_303
timestamp 1649977179
transform 1 0 28980 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_311
timestamp 1649977179
transform 1 0 29716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_323
timestamp 1649977179
transform 1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1649977179
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_341
timestamp 1649977179
transform 1 0 32476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_353
timestamp 1649977179
transform 1 0 33580 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_359
timestamp 1649977179
transform 1 0 34132 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_367
timestamp 1649977179
transform 1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_425
timestamp 1649977179
transform 1 0 40204 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_431
timestamp 1649977179
transform 1 0 40756 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_438
timestamp 1649977179
transform 1 0 41400 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_446
timestamp 1649977179
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_488
timestamp 1649977179
transform 1 0 46000 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_495
timestamp 1649977179
transform 1 0 46644 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_508
timestamp 1649977179
transform 1 0 47840 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1649977179
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_207
timestamp 1649977179
transform 1 0 20148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_219
timestamp 1649977179
transform 1 0 21252 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_230
timestamp 1649977179
transform 1 0 22264 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_241
timestamp 1649977179
transform 1 0 23276 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1649977179
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_263
timestamp 1649977179
transform 1 0 25300 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_269
timestamp 1649977179
transform 1 0 25852 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_278
timestamp 1649977179
transform 1 0 26680 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_284
timestamp 1649977179
transform 1 0 27232 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_353
timestamp 1649977179
transform 1 0 33580 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1649977179
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_372
timestamp 1649977179
transform 1 0 35328 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_384
timestamp 1649977179
transform 1 0 36432 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_393
timestamp 1649977179
transform 1 0 37260 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_400
timestamp 1649977179
transform 1 0 37904 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_407
timestamp 1649977179
transform 1 0 38548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_429
timestamp 1649977179
transform 1 0 40572 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_436
timestamp 1649977179
transform 1 0 41216 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_448
timestamp 1649977179
transform 1 0 42320 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_456
timestamp 1649977179
transform 1 0 43056 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_462
timestamp 1649977179
transform 1 0 43608 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1649977179
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_177
timestamp 1649977179
transform 1 0 17388 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_189
timestamp 1649977179
transform 1 0 18492 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_201
timestamp 1649977179
transform 1 0 19596 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_213
timestamp 1649977179
transform 1 0 20700 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1649977179
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_233
timestamp 1649977179
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_239
timestamp 1649977179
transform 1 0 23092 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_263
timestamp 1649977179
transform 1 0 25300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1649977179
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_289
timestamp 1649977179
transform 1 0 27692 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_309
timestamp 1649977179
transform 1 0 29532 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_316
timestamp 1649977179
transform 1 0 30176 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_327
timestamp 1649977179
transform 1 0 31188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_345
timestamp 1649977179
transform 1 0 32844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_351
timestamp 1649977179
transform 1 0 33396 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_362
timestamp 1649977179
transform 1 0 34408 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1649977179
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_403
timestamp 1649977179
transform 1 0 38180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_415
timestamp 1649977179
transform 1 0 39284 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_423
timestamp 1649977179
transform 1 0 40020 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_430
timestamp 1649977179
transform 1 0 40664 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_437
timestamp 1649977179
transform 1 0 41308 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_445
timestamp 1649977179
transform 1 0 42044 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_455
timestamp 1649977179
transform 1 0 42964 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_481
timestamp 1649977179
transform 1 0 45356 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_493
timestamp 1649977179
transform 1 0 46460 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_501
timestamp 1649977179
transform 1 0 47196 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_508
timestamp 1649977179
transform 1 0 47840 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_261
timestamp 1649977179
transform 1 0 25116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_282
timestamp 1649977179
transform 1 0 27048 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_294
timestamp 1649977179
transform 1 0 28152 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1649977179
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_320
timestamp 1649977179
transform 1 0 30544 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_340
timestamp 1649977179
transform 1 0 32384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_352
timestamp 1649977179
transform 1 0 33488 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1649977179
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_371
timestamp 1649977179
transform 1 0 35236 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_379
timestamp 1649977179
transform 1 0 35972 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_397
timestamp 1649977179
transform 1 0 37628 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_414
timestamp 1649977179
transform 1 0 39192 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_429
timestamp 1649977179
transform 1 0 40572 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_441
timestamp 1649977179
transform 1 0 41676 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_449
timestamp 1649977179
transform 1 0 42412 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_454
timestamp 1649977179
transform 1 0 42872 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_462
timestamp 1649977179
transform 1 0 43608 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1649977179
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_309
timestamp 1649977179
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_321
timestamp 1649977179
transform 1 0 30636 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_379
timestamp 1649977179
transform 1 0 35972 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1649977179
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_400
timestamp 1649977179
transform 1 0 37904 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_408
timestamp 1649977179
transform 1 0 38640 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_425
timestamp 1649977179
transform 1 0 40204 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_465
timestamp 1649977179
transform 1 0 43884 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_477
timestamp 1649977179
transform 1 0 44988 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_483
timestamp 1649977179
transform 1 0 45540 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_500
timestamp 1649977179
transform 1 0 47104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_508
timestamp 1649977179
transform 1 0 47840 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_259
timestamp 1649977179
transform 1 0 24932 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_271
timestamp 1649977179
transform 1 0 26036 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_283
timestamp 1649977179
transform 1 0 27140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_302
timestamp 1649977179
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_353
timestamp 1649977179
transform 1 0 33580 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1649977179
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_371
timestamp 1649977179
transform 1 0 35236 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_403
timestamp 1649977179
transform 1 0 38180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_415
timestamp 1649977179
transform 1 0 39284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_429
timestamp 1649977179
transform 1 0 40572 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_440
timestamp 1649977179
transform 1 0 41584 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_449
timestamp 1649977179
transform 1 0 42412 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_460
timestamp 1649977179
transform 1 0 43424 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_472
timestamp 1649977179
transform 1 0 44528 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_482
timestamp 1649977179
transform 1 0 45448 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_492
timestamp 1649977179
transform 1 0 46368 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_512
timestamp 1649977179
transform 1 0 48208 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_245
timestamp 1649977179
transform 1 0 23644 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_252
timestamp 1649977179
transform 1 0 24288 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1649977179
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_308
timestamp 1649977179
transform 1 0 29440 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_319
timestamp 1649977179
transform 1 0 30452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_331
timestamp 1649977179
transform 1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_368
timestamp 1649977179
transform 1 0 34960 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_380
timestamp 1649977179
transform 1 0 36064 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1649977179
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_413
timestamp 1649977179
transform 1 0 39100 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_425
timestamp 1649977179
transform 1 0 40204 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_444
timestamp 1649977179
transform 1 0 41952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_453
timestamp 1649977179
transform 1 0 42780 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_460
timestamp 1649977179
transform 1 0 43424 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_480
timestamp 1649977179
transform 1 0 45264 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_489
timestamp 1649977179
transform 1 0 46092 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_500
timestamp 1649977179
transform 1 0 47104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_510
timestamp 1649977179
transform 1 0 48024 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_11
timestamp 1649977179
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_17
timestamp 1649977179
transform 1 0 2668 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_25
timestamp 1649977179
transform 1 0 3404 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_272
timestamp 1649977179
transform 1 0 26128 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_284
timestamp 1649977179
transform 1 0 27232 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_293
timestamp 1649977179
transform 1 0 28060 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1649977179
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_315
timestamp 1649977179
transform 1 0 30084 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_325
timestamp 1649977179
transform 1 0 31004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_343
timestamp 1649977179
transform 1 0 32660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_351
timestamp 1649977179
transform 1 0 33396 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1649977179
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_373
timestamp 1649977179
transform 1 0 35420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_382
timestamp 1649977179
transform 1 0 36248 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_392
timestamp 1649977179
transform 1 0 37168 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_402
timestamp 1649977179
transform 1 0 38088 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_411
timestamp 1649977179
transform 1 0 38916 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_428
timestamp 1649977179
transform 1 0 40480 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_439
timestamp 1649977179
transform 1 0 41492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_449
timestamp 1649977179
transform 1 0 42412 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_456
timestamp 1649977179
transform 1 0 43056 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1649977179
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_32
timestamp 1649977179
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_44
timestamp 1649977179
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_264
timestamp 1649977179
transform 1 0 25392 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1649977179
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_297
timestamp 1649977179
transform 1 0 28428 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_306
timestamp 1649977179
transform 1 0 29256 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_313
timestamp 1649977179
transform 1 0 29900 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_321
timestamp 1649977179
transform 1 0 30636 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_326
timestamp 1649977179
transform 1 0 31096 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1649977179
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_342
timestamp 1649977179
transform 1 0 32568 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_354
timestamp 1649977179
transform 1 0 33672 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_366
timestamp 1649977179
transform 1 0 34776 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_377
timestamp 1649977179
transform 1 0 35788 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_388
timestamp 1649977179
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_401
timestamp 1649977179
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_410
timestamp 1649977179
transform 1 0 38824 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_420
timestamp 1649977179
transform 1 0 39744 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_427
timestamp 1649977179
transform 1 0 40388 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_434
timestamp 1649977179
transform 1 0 41032 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_452
timestamp 1649977179
transform 1 0 42688 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_458
timestamp 1649977179
transform 1 0 43240 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_464
timestamp 1649977179
transform 1 0 43792 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_471
timestamp 1649977179
transform 1 0 44436 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_483
timestamp 1649977179
transform 1 0 45540 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_495
timestamp 1649977179
transform 1 0 46644 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_508
timestamp 1649977179
transform 1 0 47840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_14
timestamp 1649977179
transform 1 0 2392 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 1649977179
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_259
timestamp 1649977179
transform 1 0 24932 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_268
timestamp 1649977179
transform 1 0 25760 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_275
timestamp 1649977179
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_287
timestamp 1649977179
transform 1 0 27508 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1649977179
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_313
timestamp 1649977179
transform 1 0 29900 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_319
timestamp 1649977179
transform 1 0 30452 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_325
timestamp 1649977179
transform 1 0 31004 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_343
timestamp 1649977179
transform 1 0 32660 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_353
timestamp 1649977179
transform 1 0 33580 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_361
timestamp 1649977179
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_385
timestamp 1649977179
transform 1 0 36524 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_395
timestamp 1649977179
transform 1 0 37444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_407
timestamp 1649977179
transform 1 0 38548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_425
timestamp 1649977179
transform 1 0 40204 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_434
timestamp 1649977179
transform 1 0 41032 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_460
timestamp 1649977179
transform 1 0 43424 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_467
timestamp 1649977179
transform 1 0 44068 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_493
timestamp 1649977179
transform 1 0 46460 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_502
timestamp 1649977179
transform 1 0 47288 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_509
timestamp 1649977179
transform 1 0 47932 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_515
timestamp 1649977179
transform 1 0 48484 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_266
timestamp 1649977179
transform 1 0 25576 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_319
timestamp 1649977179
transform 1 0 30452 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_327
timestamp 1649977179
transform 1 0 31188 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_344
timestamp 1649977179
transform 1 0 32752 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_348
timestamp 1649977179
transform 1 0 33120 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_357
timestamp 1649977179
transform 1 0 33948 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_367
timestamp 1649977179
transform 1 0 34868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_379
timestamp 1649977179
transform 1 0 35972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_435
timestamp 1649977179
transform 1 0 41124 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_439
timestamp 1649977179
transform 1 0 41492 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_469
timestamp 1649977179
transform 1 0 44252 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_476
timestamp 1649977179
transform 1 0 44896 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_488
timestamp 1649977179
transform 1 0 46000 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_496
timestamp 1649977179
transform 1 0 46736 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_500
timestamp 1649977179
transform 1 0 47104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_508
timestamp 1649977179
transform 1 0 47840 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_11
timestamp 1649977179
transform 1 0 2116 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_16
timestamp 1649977179
transform 1 0 2576 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1649977179
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_260
timestamp 1649977179
transform 1 0 25024 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_268
timestamp 1649977179
transform 1 0 25760 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_291
timestamp 1649977179
transform 1 0 27876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_303
timestamp 1649977179
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_312
timestamp 1649977179
transform 1 0 29808 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_320
timestamp 1649977179
transform 1 0 30544 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_324
timestamp 1649977179
transform 1 0 30912 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_332
timestamp 1649977179
transform 1 0 31648 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_336
timestamp 1649977179
transform 1 0 32016 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_344
timestamp 1649977179
transform 1 0 32752 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_351
timestamp 1649977179
transform 1 0 33396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_355
timestamp 1649977179
transform 1 0 33764 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1649977179
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_370
timestamp 1649977179
transform 1 0 35144 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_378
timestamp 1649977179
transform 1 0 35880 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_388
timestamp 1649977179
transform 1 0 36800 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_400
timestamp 1649977179
transform 1 0 37904 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_412
timestamp 1649977179
transform 1 0 39008 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_429
timestamp 1649977179
transform 1 0 40572 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_435
timestamp 1649977179
transform 1 0 41124 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_460
timestamp 1649977179
transform 1 0 43424 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_467
timestamp 1649977179
transform 1 0 44068 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_480
timestamp 1649977179
transform 1 0 45264 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_492
timestamp 1649977179
transform 1 0 46368 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1649977179
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_9
timestamp 1649977179
transform 1 0 1932 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_31
timestamp 1649977179
transform 1 0 3956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_43
timestamp 1649977179
transform 1 0 5060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_269
timestamp 1649977179
transform 1 0 25852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1649977179
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_287
timestamp 1649977179
transform 1 0 27508 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_307
timestamp 1649977179
transform 1 0 29348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_327
timestamp 1649977179
transform 1 0 31188 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_346
timestamp 1649977179
transform 1 0 32936 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_350
timestamp 1649977179
transform 1 0 33304 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_354
timestamp 1649977179
transform 1 0 33672 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_364
timestamp 1649977179
transform 1 0 34592 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_371
timestamp 1649977179
transform 1 0 35236 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_378
timestamp 1649977179
transform 1 0 35880 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1649977179
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_397
timestamp 1649977179
transform 1 0 37628 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_409
timestamp 1649977179
transform 1 0 38732 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_438
timestamp 1649977179
transform 1 0 41400 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_446
timestamp 1649977179
transform 1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_465
timestamp 1649977179
transform 1 0 43884 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_482
timestamp 1649977179
transform 1 0 45448 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_490
timestamp 1649977179
transform 1 0 46184 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_498
timestamp 1649977179
transform 1 0 46920 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1649977179
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_14
timestamp 1649977179
transform 1 0 2392 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1649977179
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_257
timestamp 1649977179
transform 1 0 24748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_263
timestamp 1649977179
transform 1 0 25300 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_276
timestamp 1649977179
transform 1 0 26496 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_284
timestamp 1649977179
transform 1 0 27232 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_295
timestamp 1649977179
transform 1 0 28244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_340
timestamp 1649977179
transform 1 0 32384 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_352
timestamp 1649977179
transform 1 0 33488 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_368
timestamp 1649977179
transform 1 0 34960 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_376
timestamp 1649977179
transform 1 0 35696 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_382
timestamp 1649977179
transform 1 0 36248 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_402
timestamp 1649977179
transform 1 0 38088 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_408
timestamp 1649977179
transform 1 0 38640 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_416
timestamp 1649977179
transform 1 0 39376 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_437
timestamp 1649977179
transform 1 0 41308 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_449
timestamp 1649977179
transform 1 0 42412 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_461
timestamp 1649977179
transform 1 0 43516 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_482
timestamp 1649977179
transform 1 0 45448 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_488
timestamp 1649977179
transform 1 0 46000 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_492
timestamp 1649977179
transform 1 0 46368 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1649977179
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_254
timestamp 1649977179
transform 1 0 24472 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_263
timestamp 1649977179
transform 1 0 25300 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_287
timestamp 1649977179
transform 1 0 27508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_299
timestamp 1649977179
transform 1 0 28612 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_310
timestamp 1649977179
transform 1 0 29624 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_322
timestamp 1649977179
transform 1 0 30728 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1649977179
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_344
timestamp 1649977179
transform 1 0 32752 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_356
timestamp 1649977179
transform 1 0 33856 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_368
timestamp 1649977179
transform 1 0 34960 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_378
timestamp 1649977179
transform 1 0 35880 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1649977179
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_415
timestamp 1649977179
transform 1 0 39284 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_423
timestamp 1649977179
transform 1 0 40020 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_433
timestamp 1649977179
transform 1 0 40940 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_445
timestamp 1649977179
transform 1 0 42044 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_456
timestamp 1649977179
transform 1 0 43056 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_468
timestamp 1649977179
transform 1 0 44160 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_478
timestamp 1649977179
transform 1 0 45080 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_488
timestamp 1649977179
transform 1 0 46000 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_498
timestamp 1649977179
transform 1 0 46920 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_510
timestamp 1649977179
transform 1 0 48024 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_212
timestamp 1649977179
transform 1 0 20608 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_224
timestamp 1649977179
transform 1 0 21712 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_236
timestamp 1649977179
transform 1 0 22816 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1649977179
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_269
timestamp 1649977179
transform 1 0 25852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_286
timestamp 1649977179
transform 1 0 27416 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1649977179
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1649977179
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_314
timestamp 1649977179
transform 1 0 29992 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_326
timestamp 1649977179
transform 1 0 31096 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_338
timestamp 1649977179
transform 1 0 32200 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_350
timestamp 1649977179
transform 1 0 33304 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1649977179
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_375
timestamp 1649977179
transform 1 0 35604 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_386
timestamp 1649977179
transform 1 0 36616 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_398
timestamp 1649977179
transform 1 0 37720 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_410
timestamp 1649977179
transform 1 0 38824 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_418
timestamp 1649977179
transform 1 0 39560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_428
timestamp 1649977179
transform 1 0 40480 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_448
timestamp 1649977179
transform 1 0 42320 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_468
timestamp 1649977179
transform 1 0 44160 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_492
timestamp 1649977179
transform 1 0 46368 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_512
timestamp 1649977179
transform 1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_265
timestamp 1649977179
transform 1 0 25484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1649977179
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_297
timestamp 1649977179
transform 1 0 28428 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_365
timestamp 1649977179
transform 1 0 34684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_383
timestamp 1649977179
transform 1 0 36340 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_411
timestamp 1649977179
transform 1 0 38916 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_432
timestamp 1649977179
transform 1 0 40848 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_439
timestamp 1649977179
transform 1 0 41492 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_479
timestamp 1649977179
transform 1 0 45172 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_491
timestamp 1649977179
transform 1 0 46276 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_500
timestamp 1649977179
transform 1 0 47104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_508
timestamp 1649977179
transform 1 0 47840 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_260
timestamp 1649977179
transform 1 0 25024 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1649977179
transform 1 0 26220 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_284
timestamp 1649977179
transform 1 0 27232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_291
timestamp 1649977179
transform 1 0 27876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_295
timestamp 1649977179
transform 1 0 28244 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1649977179
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_313
timestamp 1649977179
transform 1 0 29900 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_325
timestamp 1649977179
transform 1 0 31004 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_337
timestamp 1649977179
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_349
timestamp 1649977179
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1649977179
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1649977179
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_380
timestamp 1649977179
transform 1 0 36064 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_390
timestamp 1649977179
transform 1 0 36984 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_402
timestamp 1649977179
transform 1 0 38088 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_414
timestamp 1649977179
transform 1 0 39192 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_426
timestamp 1649977179
transform 1 0 40296 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_435
timestamp 1649977179
transform 1 0 41124 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_442
timestamp 1649977179
transform 1 0 41768 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_454
timestamp 1649977179
transform 1 0 42872 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_462
timestamp 1649977179
transform 1 0 43608 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_470
timestamp 1649977179
transform 1 0 44344 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1649977179
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_257
timestamp 1649977179
transform 1 0 24748 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1649977179
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_321
timestamp 1649977179
transform 1 0 30636 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_331
timestamp 1649977179
transform 1 0 31556 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_353
timestamp 1649977179
transform 1 0 33580 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_365
timestamp 1649977179
transform 1 0 34684 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_371
timestamp 1649977179
transform 1 0 35236 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_380
timestamp 1649977179
transform 1 0 36064 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_387
timestamp 1649977179
transform 1 0 36708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_409
timestamp 1649977179
transform 1 0 38732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_434
timestamp 1649977179
transform 1 0 41032 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_443
timestamp 1649977179
transform 1 0 41860 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_468
timestamp 1649977179
transform 1 0 44160 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_480
timestamp 1649977179
transform 1 0 45264 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_500
timestamp 1649977179
transform 1 0 47104 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_508
timestamp 1649977179
transform 1 0 47840 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_269
timestamp 1649977179
transform 1 0 25852 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_281
timestamp 1649977179
transform 1 0 26956 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_293
timestamp 1649977179
transform 1 0 28060 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_297
timestamp 1649977179
transform 1 0 28428 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_303
timestamp 1649977179
transform 1 0 28980 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_319
timestamp 1649977179
transform 1 0 30452 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_339
timestamp 1649977179
transform 1 0 32292 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_346
timestamp 1649977179
transform 1 0 32936 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_358
timestamp 1649977179
transform 1 0 34040 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_66_381
timestamp 1649977179
transform 1 0 36156 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_408
timestamp 1649977179
transform 1 0 38640 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_439
timestamp 1649977179
transform 1 0 41492 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_449
timestamp 1649977179
transform 1 0 42412 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_455
timestamp 1649977179
transform 1 0 42964 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_472
timestamp 1649977179
transform 1 0 44528 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_482
timestamp 1649977179
transform 1 0 45448 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_486
timestamp 1649977179
transform 1 0 45816 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_492
timestamp 1649977179
transform 1 0 46368 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_499
timestamp 1649977179
transform 1 0 47012 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_506
timestamp 1649977179
transform 1 0 47656 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_514
timestamp 1649977179
transform 1 0 48392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_311
timestamp 1649977179
transform 1 0 29716 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_321
timestamp 1649977179
transform 1 0 30636 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_332
timestamp 1649977179
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_342
timestamp 1649977179
transform 1 0 32568 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_370
timestamp 1649977179
transform 1 0 35144 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_379
timestamp 1649977179
transform 1 0 35972 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_386
timestamp 1649977179
transform 1 0 36616 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_399
timestamp 1649977179
transform 1 0 37812 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_406
timestamp 1649977179
transform 1 0 38456 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_410
timestamp 1649977179
transform 1 0 38824 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_419
timestamp 1649977179
transform 1 0 39652 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_426
timestamp 1649977179
transform 1 0 40296 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_430
timestamp 1649977179
transform 1 0 40664 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_438
timestamp 1649977179
transform 1 0 41400 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_446
timestamp 1649977179
transform 1 0 42136 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_465
timestamp 1649977179
transform 1 0 43884 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_477
timestamp 1649977179
transform 1 0 44988 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_495
timestamp 1649977179
transform 1 0 46644 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_508
timestamp 1649977179
transform 1 0 47840 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_269
timestamp 1649977179
transform 1 0 25852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_278
timestamp 1649977179
transform 1 0 26680 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_286
timestamp 1649977179
transform 1 0 27416 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_295
timestamp 1649977179
transform 1 0 28244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_302
timestamp 1649977179
transform 1 0 28888 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_326
timestamp 1649977179
transform 1 0 31096 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_339
timestamp 1649977179
transform 1 0 32292 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_344
timestamp 1649977179
transform 1 0 32752 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_356
timestamp 1649977179
transform 1 0 33856 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_374
timestamp 1649977179
transform 1 0 35512 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_386
timestamp 1649977179
transform 1 0 36616 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_398
timestamp 1649977179
transform 1 0 37720 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_410
timestamp 1649977179
transform 1 0 38824 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_418
timestamp 1649977179
transform 1 0 39560 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_68_446
timestamp 1649977179
transform 1 0 42136 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_452
timestamp 1649977179
transform 1 0 42688 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_456
timestamp 1649977179
transform 1 0 43056 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_468
timestamp 1649977179
transform 1 0 44160 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1649977179
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_69_248
timestamp 1649977179
transform 1 0 23920 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_69_270
timestamp 1649977179
transform 1 0 25944 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_278
timestamp 1649977179
transform 1 0 26680 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_299
timestamp 1649977179
transform 1 0 28612 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_306
timestamp 1649977179
transform 1 0 29256 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_468
timestamp 1649977179
transform 1 0 44160 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_476
timestamp 1649977179
transform 1 0 44896 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_493
timestamp 1649977179
transform 1 0 46460 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_500
timestamp 1649977179
transform 1 0 47104 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1649977179
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_88
timestamp 1649977179
transform 1 0 9200 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_100
timestamp 1649977179
transform 1 0 10304 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_112
timestamp 1649977179
transform 1 0 11408 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_124
timestamp 1649977179
transform 1 0 12512 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_136
timestamp 1649977179
transform 1 0 13616 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_237
timestamp 1649977179
transform 1 0 22908 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_244
timestamp 1649977179
transform 1 0 23552 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_256
timestamp 1649977179
transform 1 0 24656 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_276
timestamp 1649977179
transform 1 0 26496 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_285
timestamp 1649977179
transform 1 0 27324 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_295
timestamp 1649977179
transform 1 0 28244 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1649977179
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_325
timestamp 1649977179
transform 1 0 31004 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_337
timestamp 1649977179
transform 1 0 32108 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_349
timestamp 1649977179
transform 1 0 33212 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_356
timestamp 1649977179
transform 1 0 33856 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_373
timestamp 1649977179
transform 1 0 35420 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_381
timestamp 1649977179
transform 1 0 36156 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_386
timestamp 1649977179
transform 1 0 36616 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_397
timestamp 1649977179
transform 1 0 37628 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_406
timestamp 1649977179
transform 1 0 38456 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_441
timestamp 1649977179
transform 1 0 41676 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_451
timestamp 1649977179
transform 1 0 42596 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_460
timestamp 1649977179
transform 1 0 43424 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_512
timestamp 1649977179
transform 1 0 48208 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_175
timestamp 1649977179
transform 1 0 17204 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_187
timestamp 1649977179
transform 1 0 18308 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_199
timestamp 1649977179
transform 1 0 19412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_211
timestamp 1649977179
transform 1 0 20516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_266
timestamp 1649977179
transform 1 0 25576 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_275
timestamp 1649977179
transform 1 0 26404 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_310
timestamp 1649977179
transform 1 0 29624 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_322
timestamp 1649977179
transform 1 0 30728 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_328
timestamp 1649977179
transform 1 0 31280 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_356
timestamp 1649977179
transform 1 0 33856 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_367
timestamp 1649977179
transform 1 0 34868 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_377
timestamp 1649977179
transform 1 0 35788 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_381
timestamp 1649977179
transform 1 0 36156 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_388
timestamp 1649977179
transform 1 0 36800 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_397
timestamp 1649977179
transform 1 0 37628 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_437
timestamp 1649977179
transform 1 0 41308 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_444
timestamp 1649977179
transform 1 0 41952 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_456
timestamp 1649977179
transform 1 0 43056 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_464
timestamp 1649977179
transform 1 0 43792 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_482
timestamp 1649977179
transform 1 0 45448 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_489
timestamp 1649977179
transform 1 0 46092 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_500
timestamp 1649977179
transform 1 0 47104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_508
timestamp 1649977179
transform 1 0 47840 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_273
timestamp 1649977179
transform 1 0 26220 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_292
timestamp 1649977179
transform 1 0 27968 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1649977179
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_325
timestamp 1649977179
transform 1 0 31004 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_354
timestamp 1649977179
transform 1 0 33672 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_362
timestamp 1649977179
transform 1 0 34408 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_387
timestamp 1649977179
transform 1 0 36708 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_407
timestamp 1649977179
transform 1 0 38548 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_416
timestamp 1649977179
transform 1 0 39376 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_426
timestamp 1649977179
transform 1 0 40296 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_434
timestamp 1649977179
transform 1 0 41032 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_451
timestamp 1649977179
transform 1 0 42596 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_471
timestamp 1649977179
transform 1 0 44436 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_483
timestamp 1649977179
transform 1 0 45540 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1649977179
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_284
timestamp 1649977179
transform 1 0 27232 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_299
timestamp 1649977179
transform 1 0 28612 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_311
timestamp 1649977179
transform 1 0 29716 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_323
timestamp 1649977179
transform 1 0 30820 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_330
timestamp 1649977179
transform 1 0 31464 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_344
timestamp 1649977179
transform 1 0 32752 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_364
timestamp 1649977179
transform 1 0 34592 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_380
timestamp 1649977179
transform 1 0 36064 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_387
timestamp 1649977179
transform 1 0 36708 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_398
timestamp 1649977179
transform 1 0 37720 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_410
timestamp 1649977179
transform 1 0 38824 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_422
timestamp 1649977179
transform 1 0 39928 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_428
timestamp 1649977179
transform 1 0 40480 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_436
timestamp 1649977179
transform 1 0 41216 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_444
timestamp 1649977179
transform 1 0 41952 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_454
timestamp 1649977179
transform 1 0 42872 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_500
timestamp 1649977179
transform 1 0 47104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_508
timestamp 1649977179
transform 1 0 47840 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_32
timestamp 1649977179
transform 1 0 4048 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_44
timestamp 1649977179
transform 1 0 5152 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_56
timestamp 1649977179
transform 1 0 6256 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_68
timestamp 1649977179
transform 1 0 7360 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1649977179
transform 1 0 8464 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_286
timestamp 1649977179
transform 1 0 27416 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_290
timestamp 1649977179
transform 1 0 27784 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_297
timestamp 1649977179
transform 1 0 28428 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_305
timestamp 1649977179
transform 1 0 29164 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_351
timestamp 1649977179
transform 1 0 33396 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_355
timestamp 1649977179
transform 1 0 33764 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_480
timestamp 1649977179
transform 1 0 45264 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_487
timestamp 1649977179
transform 1 0 45908 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1649977179
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_32
timestamp 1649977179
transform 1 0 4048 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_44
timestamp 1649977179
transform 1 0 5152 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_444
timestamp 1649977179
transform 1 0 41952 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_489
timestamp 1649977179
transform 1 0 46092 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_496
timestamp 1649977179
transform 1 0 46736 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_508
timestamp 1649977179
transform 1 0 47840 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_14
timestamp 1649977179
transform 1 0 2392 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_26
timestamp 1649977179
transform 1 0 3496 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_428
timestamp 1649977179
transform 1 0 40480 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_440
timestamp 1649977179
transform 1 0 41584 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_452
timestamp 1649977179
transform 1 0 42688 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_464
timestamp 1649977179
transform 1 0 43792 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1649977179
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_85
timestamp 1649977179
transform 1 0 8924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_95
timestamp 1649977179
transform 1 0 9844 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_107
timestamp 1649977179
transform 1 0 10948 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_489
timestamp 1649977179
transform 1 0 46092 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1649977179
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1649977179
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1649977179
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_10
timestamp 1649977179
transform 1 0 2024 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_17
timestamp 1649977179
transform 1 0 2668 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_24
timestamp 1649977179
transform 1 0 3312 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_32
timestamp 1649977179
transform 1 0 4048 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_44
timestamp 1649977179
transform 1 0 5152 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_56
timestamp 1649977179
transform 1 0 6256 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_68
timestamp 1649977179
transform 1 0 7360 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_80
timestamp 1649977179
transform 1 0 8464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_96
timestamp 1649977179
transform 1 0 9936 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_108
timestamp 1649977179
transform 1 0 11040 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_120
timestamp 1649977179
transform 1 0 12144 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_132
timestamp 1649977179
transform 1 0 13248 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_281
timestamp 1649977179
transform 1 0 26956 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_288
timestamp 1649977179
transform 1 0 27600 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_300
timestamp 1649977179
transform 1 0 28704 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_316
timestamp 1649977179
transform 1 0 30176 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_328
timestamp 1649977179
transform 1 0 31280 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_340
timestamp 1649977179
transform 1 0 32384 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_352
timestamp 1649977179
transform 1 0 33488 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_405
timestamp 1649977179
transform 1 0 38364 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_417
timestamp 1649977179
transform 1 0 39468 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_444
timestamp 1649977179
transform 1 0 41952 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_456
timestamp 1649977179
transform 1 0 43056 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_468
timestamp 1649977179
transform 1 0 44160 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_483
timestamp 1649977179
transform 1 0 45540 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1649977179
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1649977179
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_9
timestamp 1649977179
transform 1 0 1932 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_34
timestamp 1649977179
transform 1 0 4232 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_46
timestamp 1649977179
transform 1 0 5336 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_50
timestamp 1649977179
transform 1 0 5704 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_77
timestamp 1649977179
transform 1 0 8188 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_82
timestamp 1649977179
transform 1 0 8648 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_95
timestamp 1649977179
transform 1 0 9844 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_108
timestamp 1649977179
transform 1 0 11040 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_116
timestamp 1649977179
transform 1 0 11776 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_127
timestamp 1649977179
transform 1 0 12788 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_152
timestamp 1649977179
transform 1 0 15088 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_156
timestamp 1649977179
transform 1 0 15456 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_160
timestamp 1649977179
transform 1 0 15824 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_233
timestamp 1649977179
transform 1 0 22540 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_239
timestamp 1649977179
transform 1 0 23092 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_251
timestamp 1649977179
transform 1 0 24196 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_258
timestamp 1649977179
transform 1 0 24840 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_265
timestamp 1649977179
transform 1 0 25484 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_79_274
timestamp 1649977179
transform 1 0 26312 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_285
timestamp 1649977179
transform 1 0 27324 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_297
timestamp 1649977179
transform 1 0 28428 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_320
timestamp 1649977179
transform 1 0 30544 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_332
timestamp 1649977179
transform 1 0 31648 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_377
timestamp 1649977179
transform 1 0 35788 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_381
timestamp 1649977179
transform 1 0 36156 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_389
timestamp 1649977179
transform 1 0 36892 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_401
timestamp 1649977179
transform 1 0 37996 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_423
timestamp 1649977179
transform 1 0 40020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_435
timestamp 1649977179
transform 1 0 41124 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1649977179
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1649977179
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1649977179
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_35
timestamp 1649977179
transform 1 0 4324 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_43
timestamp 1649977179
transform 1 0 5060 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_66
timestamp 1649977179
transform 1 0 7176 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_78
timestamp 1649977179
transform 1 0 8280 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_96
timestamp 1649977179
transform 1 0 9936 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_104
timestamp 1649977179
transform 1 0 10672 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_127
timestamp 1649977179
transform 1 0 12788 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_134
timestamp 1649977179
transform 1 0 13432 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_147
timestamp 1649977179
transform 1 0 14628 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_176
timestamp 1649977179
transform 1 0 17296 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_188
timestamp 1649977179
transform 1 0 18400 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_239
timestamp 1649977179
transform 1 0 23092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_302
timestamp 1649977179
transform 1 0 28888 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_312
timestamp 1649977179
transform 1 0 29808 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_324
timestamp 1649977179
transform 1 0 30912 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_336
timestamp 1649977179
transform 1 0 32016 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_347
timestamp 1649977179
transform 1 0 33028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_359
timestamp 1649977179
transform 1 0 34132 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_373
timestamp 1649977179
transform 1 0 35420 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_397
timestamp 1649977179
transform 1 0 37628 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_405
timestamp 1649977179
transform 1 0 38364 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_417
timestamp 1649977179
transform 1 0 39468 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_439
timestamp 1649977179
transform 1 0 41492 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_461
timestamp 1649977179
transform 1 0 43516 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_473
timestamp 1649977179
transform 1 0 44620 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_483
timestamp 1649977179
transform 1 0 45540 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1649977179
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1649977179
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1649977179
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1649977179
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_138
timestamp 1649977179
transform 1 0 13800 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_163
timestamp 1649977179
transform 1 0 16100 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_229
timestamp 1649977179
transform 1 0 22172 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_251
timestamp 1649977179
transform 1 0 24196 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_276
timestamp 1649977179
transform 1 0 26496 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_302
timestamp 1649977179
transform 1 0 28888 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_310
timestamp 1649977179
transform 1 0 29624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1649977179
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_343
timestamp 1649977179
transform 1 0 32660 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_365
timestamp 1649977179
transform 1 0 34684 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_380
timestamp 1649977179
transform 1 0 36064 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_387
timestamp 1649977179
transform 1 0 36708 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_414
timestamp 1649977179
transform 1 0 39192 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_426
timestamp 1649977179
transform 1 0 40296 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_438
timestamp 1649977179
transform 1 0 41400 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_443
timestamp 1649977179
transform 1 0 41860 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1649977179
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_508
timestamp 1649977179
transform 1 0 47840 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1649977179
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_17
timestamp 1649977179
transform 1 0 2668 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1649977179
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_35
timestamp 1649977179
transform 1 0 4324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_42
timestamp 1649977179
transform 1 0 4968 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_49
timestamp 1649977179
transform 1 0 5612 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_55
timestamp 1649977179
transform 1 0 6164 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_57
timestamp 1649977179
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_69
timestamp 1649977179
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1649977179
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_88
timestamp 1649977179
transform 1 0 9200 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_100
timestamp 1649977179
transform 1 0 10304 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_113
timestamp 1649977179
transform 1 0 11500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_127
timestamp 1649977179
transform 1 0 12788 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_131
timestamp 1649977179
transform 1 0 13156 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1649977179
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_146
timestamp 1649977179
transform 1 0 14536 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_154
timestamp 1649977179
transform 1 0 15272 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_82_159
timestamp 1649977179
transform 1 0 15732 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_167
timestamp 1649977179
transform 1 0 16468 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_169
timestamp 1649977179
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_181
timestamp 1649977179
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1649977179
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_225
timestamp 1649977179
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_237
timestamp 1649977179
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1649977179
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_259
timestamp 1649977179
transform 1 0 24932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_266
timestamp 1649977179
transform 1 0 25576 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_272
timestamp 1649977179
transform 1 0 26128 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_276
timestamp 1649977179
transform 1 0 26496 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_281
timestamp 1649977179
transform 1 0 26956 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_293
timestamp 1649977179
transform 1 0 28060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1649977179
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_316
timestamp 1649977179
transform 1 0 30176 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_328
timestamp 1649977179
transform 1 0 31280 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_337
timestamp 1649977179
transform 1 0 32108 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_348
timestamp 1649977179
transform 1 0 33120 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_360
timestamp 1649977179
transform 1 0 34224 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_381
timestamp 1649977179
transform 1 0 36156 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_393
timestamp 1649977179
transform 1 0 37260 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_405
timestamp 1649977179
transform 1 0 38364 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_417
timestamp 1649977179
transform 1 0 39468 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_449
timestamp 1649977179
transform 1 0 42412 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_461
timestamp 1649977179
transform 1 0 43516 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_473
timestamp 1649977179
transform 1 0 44620 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_493
timestamp 1649977179
transform 1 0 46460 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_500
timestamp 1649977179
transform 1 0 47104 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_508
timestamp 1649977179
transform 1 0 47840 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0708_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16928 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0710_
timestamp 1649977179
transform 1 0 19596 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0711_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19780 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1649977179
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1649977179
transform 1 0 46460 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0722_
timestamp 1649977179
transform 1 0 8280 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0723_
timestamp 1649977179
transform 1 0 10212 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1649977179
transform 1 0 26036 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1649977179
transform 1 0 4048 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1649977179
transform 1 0 47380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0729_
timestamp 1649977179
transform 1 0 9108 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1649977179
transform 1 0 5428 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1649977179
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0735_
timestamp 1649977179
transform 1 0 9016 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1649977179
transform 1 0 29900 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1649977179
transform 1 0 1472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0741_
timestamp 1649977179
transform 1 0 9016 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1649977179
transform 1 0 32752 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1649977179
transform 1 0 47564 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1649977179
transform 1 0 46184 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0747_
timestamp 1649977179
transform 1 0 9108 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1649977179
transform 1 0 46368 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1649977179
transform 1 0 22816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0753_
timestamp 1649977179
transform 1 0 15824 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  _0754_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16560 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1649977179
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1649977179
transform 1 0 45264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1649977179
transform 1 0 45908 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1649977179
transform 1 0 2300 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0766_
timestamp 1649977179
transform 1 0 18032 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1649977179
transform 1 0 40204 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1649977179
transform 1 0 21988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1649977179
transform 1 0 16928 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1649977179
transform 1 0 41124 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0772_
timestamp 1649977179
transform 1 0 16836 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1649977179
transform 1 0 32200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1649977179
transform 1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1649977179
transform 1 0 35880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0778_
timestamp 1649977179
transform 1 0 17940 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1649977179
transform 1 0 38088 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1649977179
transform 1 0 45632 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0784_
timestamp 1649977179
transform 1 0 7728 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0785_
timestamp 1649977179
transform 1 0 9108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1649977179
transform 1 0 15548 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1649977179
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1649977179
transform 1 0 3036 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1649977179
transform 1 0 38640 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0791_
timestamp 1649977179
transform 1 0 7912 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1649977179
transform 1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1649977179
transform 1 0 41676 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1649977179
transform 1 0 25392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1649977179
transform 1 0 2392 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0797_
timestamp 1649977179
transform 1 0 7820 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1649977179
transform 1 0 13064 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1649977179
transform 1 0 12512 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1649977179
transform 1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1649977179
transform 1 0 13156 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0803_
timestamp 1649977179
transform 1 0 7820 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1649977179
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1649977179
transform 1 0 46184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0809_
timestamp 1649977179
transform 1 0 7452 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1649977179
transform 1 0 35788 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1649977179
transform 1 0 14352 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0815_
timestamp 1649977179
transform 1 0 17664 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1649977179
transform 1 0 24564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1649977179
transform 1 0 25208 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0821_
timestamp 1649977179
transform 1 0 17756 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1649977179
transform 1 0 2576 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1649977179
transform 1 0 40756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1649977179
transform 1 0 41676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1649977179
transform 1 0 2760 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0827_
timestamp 1649977179
transform 1 0 16836 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1649977179
transform 1 0 2300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1649977179
transform 1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1649977179
transform 1 0 2760 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0833_
timestamp 1649977179
transform 1 0 17664 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1649977179
transform 1 0 46736 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1649977179
transform 1 0 2300 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1649977179
transform 1 0 40020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1649977179
transform 1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1649977179
transform 1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1649977179
transform 1 0 27324 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1649977179
transform 1 0 26404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1649977179
transform 1 0 26680 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1649977179
transform 1 0 37904 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1649977179
transform 1 0 37720 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1649977179
transform 1 0 38640 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0846_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0847_
timestamp 1649977179
transform 1 0 46184 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1649977179
transform 1 0 35604 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1649977179
transform 1 0 34408 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0850_
timestamp 1649977179
transform 1 0 46184 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1649977179
transform 1 0 35604 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0852_
timestamp 1649977179
transform 1 0 37904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1649977179
transform 1 0 39100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37444 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38272 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38916 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0860_
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0861_
timestamp 1649977179
transform 1 0 39928 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0862_
timestamp 1649977179
transform 1 0 40296 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0863_
timestamp 1649977179
transform 1 0 39284 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1649977179
transform 1 0 42780 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0865_
timestamp 1649977179
transform 1 0 43240 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42780 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0867_
timestamp 1649977179
transform 1 0 41308 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0868_
timestamp 1649977179
transform 1 0 40572 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1649977179
transform 1 0 24748 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1649977179
transform 1 0 21988 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1649977179
transform 1 0 26680 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1649977179
transform 1 0 27876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1649977179
transform 1 0 27600 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0876_
timestamp 1649977179
transform 1 0 31004 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1649977179
transform 1 0 30360 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1649977179
transform 1 0 31004 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31280 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0880_
timestamp 1649977179
transform 1 0 30820 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0881_
timestamp 1649977179
transform 1 0 28336 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0882_
timestamp 1649977179
transform 1 0 27232 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0883_
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0884_
timestamp 1649977179
transform 1 0 25392 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0885_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0886_
timestamp 1649977179
transform 1 0 36156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _0887_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23920 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0888_
timestamp 1649977179
transform 1 0 41400 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0889_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40112 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1649977179
transform 1 0 41032 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1649977179
transform 1 0 38272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1649977179
transform 1 0 37628 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1649977179
transform 1 0 35144 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0895_
timestamp 1649977179
transform 1 0 36156 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1649977179
transform 1 0 33856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1649977179
transform 1 0 33856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0898_
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _0899_
timestamp 1649977179
transform 1 0 33764 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33120 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1649977179
transform 1 0 34776 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0904_
timestamp 1649977179
transform 1 0 33856 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0905_
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0906_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0907_
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _0908_
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1649977179
transform 1 0 36708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0910_
timestamp 1649977179
transform 1 0 38364 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0911_
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0912_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40572 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 1649977179
transform 1 0 41216 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0914_
timestamp 1649977179
transform 1 0 35696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0915_
timestamp 1649977179
transform 1 0 32292 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0917_
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0919_
timestamp 1649977179
transform 1 0 33028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0920_
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0922_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38640 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0923_
timestamp 1649977179
transform 1 0 42504 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0924_
timestamp 1649977179
transform 1 0 30820 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0925_
timestamp 1649977179
transform 1 0 40204 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0926_
timestamp 1649977179
transform 1 0 39284 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0927_
timestamp 1649977179
transform 1 0 39836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0928_
timestamp 1649977179
transform 1 0 38456 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0929_
timestamp 1649977179
transform 1 0 37904 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0931_
timestamp 1649977179
transform 1 0 35604 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1649977179
transform 1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 35052 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0934_
timestamp 1649977179
transform 1 0 36156 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0935_
timestamp 1649977179
transform 1 0 36432 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0937_
timestamp 1649977179
transform 1 0 35880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0938_
timestamp 1649977179
transform 1 0 35880 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0940_
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0941_
timestamp 1649977179
transform 1 0 30452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0942_
timestamp 1649977179
transform 1 0 29992 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0943_
timestamp 1649977179
transform 1 0 31004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1649977179
transform 1 0 30176 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0945_
timestamp 1649977179
transform 1 0 30176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0946_
timestamp 1649977179
transform 1 0 27784 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0947_
timestamp 1649977179
transform 1 0 29348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0948_
timestamp 1649977179
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1649977179
transform 1 0 28612 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0950_
timestamp 1649977179
transform 1 0 27324 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0951_
timestamp 1649977179
transform 1 0 26864 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1649977179
transform 1 0 27048 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0953_
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0954_
timestamp 1649977179
transform 1 0 26220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0955_
timestamp 1649977179
transform 1 0 25852 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0956_
timestamp 1649977179
transform 1 0 26220 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0957_
timestamp 1649977179
transform 1 0 27048 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0958_
timestamp 1649977179
transform 1 0 25024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0959_
timestamp 1649977179
transform 1 0 24380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0960_
timestamp 1649977179
transform 1 0 24104 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0961_
timestamp 1649977179
transform 1 0 33304 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0962_
timestamp 1649977179
transform 1 0 32384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0963_
timestamp 1649977179
transform 1 0 36340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0964_
timestamp 1649977179
transform 1 0 33672 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0965_
timestamp 1649977179
transform 1 0 32752 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0966_
timestamp 1649977179
transform 1 0 40204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0967_
timestamp 1649977179
transform 1 0 32660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0968_
timestamp 1649977179
transform 1 0 33396 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0969_
timestamp 1649977179
transform 1 0 32844 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0970_
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0971_
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0972_
timestamp 1649977179
transform 1 0 35420 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0973_
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0974_
timestamp 1649977179
transform 1 0 36984 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0975_
timestamp 1649977179
transform 1 0 38272 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0976_
timestamp 1649977179
transform 1 0 38088 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0977_
timestamp 1649977179
transform 1 0 38916 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0978_
timestamp 1649977179
transform 1 0 40572 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0979_
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0980_
timestamp 1649977179
transform 1 0 41124 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0981_
timestamp 1649977179
transform 1 0 40388 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0982_
timestamp 1649977179
transform 1 0 40388 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1649977179
transform 1 0 43056 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1649977179
transform 1 0 43976 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0985_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44528 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0986_
timestamp 1649977179
transform 1 0 43608 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0987_
timestamp 1649977179
transform 1 0 45448 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0988_
timestamp 1649977179
transform 1 0 46276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0989_
timestamp 1649977179
transform 1 0 43884 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0990_
timestamp 1649977179
transform 1 0 43240 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0991_
timestamp 1649977179
transform 1 0 41584 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0992_
timestamp 1649977179
transform 1 0 39008 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0993_
timestamp 1649977179
transform 1 0 38916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0994_
timestamp 1649977179
transform 1 0 45356 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0995_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0996_
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0997_
timestamp 1649977179
transform 1 0 44160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0998_
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0999_
timestamp 1649977179
transform 1 0 43056 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1000_
timestamp 1649977179
transform 1 0 43976 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1001_
timestamp 1649977179
transform 1 0 43792 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1002_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43700 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1003_
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1004_
timestamp 1649977179
transform 1 0 40204 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1005_
timestamp 1649977179
transform 1 0 31004 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1006_
timestamp 1649977179
transform 1 0 45632 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1007_
timestamp 1649977179
transform 1 0 45172 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1649977179
transform 1 0 45264 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1011_
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44988 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1013_
timestamp 1649977179
transform 1 0 45632 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1014_
timestamp 1649977179
transform 1 0 42872 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1015_
timestamp 1649977179
transform 1 0 43976 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1016_
timestamp 1649977179
transform 1 0 42780 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1017_
timestamp 1649977179
transform 1 0 42596 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1019_
timestamp 1649977179
transform 1 0 41676 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1020_
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1021_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1022_
timestamp 1649977179
transform 1 0 45448 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1649977179
transform 1 0 44068 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1649977179
transform 1 0 44068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1025_
timestamp 1649977179
transform 1 0 44344 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1026_
timestamp 1649977179
transform 1 0 44528 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1027_
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1028_
timestamp 1649977179
transform 1 0 43148 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1029_
timestamp 1649977179
transform 1 0 42504 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 41768 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 1649977179
transform 1 0 40388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1033_
timestamp 1649977179
transform 1 0 41032 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1649977179
transform 1 0 40940 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1035_
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1036_
timestamp 1649977179
transform 1 0 43516 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1037_
timestamp 1649977179
transform 1 0 39928 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1038_
timestamp 1649977179
transform 1 0 40388 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1649977179
transform 1 0 40204 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1040_
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1041_
timestamp 1649977179
transform 1 0 37628 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1042_
timestamp 1649977179
transform 1 0 38640 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1649977179
transform 1 0 38732 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1044_
timestamp 1649977179
transform 1 0 38364 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1045_
timestamp 1649977179
transform 1 0 29992 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1046_
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1047_
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1048_
timestamp 1649977179
transform 1 0 43976 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1049_
timestamp 1649977179
transform 1 0 30452 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1050_
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 1649977179
transform 1 0 27600 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 1649977179
transform 1 0 29624 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1053_
timestamp 1649977179
transform 1 0 28244 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1054_
timestamp 1649977179
transform 1 0 27324 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1055_
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1056_
timestamp 1649977179
transform 1 0 27324 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1057_
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1058_
timestamp 1649977179
transform 1 0 31096 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1059_
timestamp 1649977179
transform 1 0 28520 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1060_
timestamp 1649977179
transform 1 0 28428 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1061_
timestamp 1649977179
transform 1 0 27324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1062_
timestamp 1649977179
transform 1 0 22908 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1063_
timestamp 1649977179
transform 1 0 29900 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1064_
timestamp 1649977179
transform 1 0 28612 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1065_
timestamp 1649977179
transform 1 0 29256 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1066_
timestamp 1649977179
transform 1 0 29900 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1067_
timestamp 1649977179
transform 1 0 30912 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1068_
timestamp 1649977179
transform 1 0 32752 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1069_
timestamp 1649977179
transform 1 0 29808 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1070_
timestamp 1649977179
transform 1 0 28520 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1071_
timestamp 1649977179
transform 1 0 28244 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1072_
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1073_
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1074_
timestamp 1649977179
transform 1 0 28244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1075_
timestamp 1649977179
transform 1 0 30728 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1076_
timestamp 1649977179
transform 1 0 28060 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1077_
timestamp 1649977179
transform 1 0 27968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1078_
timestamp 1649977179
transform 1 0 27600 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 1649977179
transform 1 0 29532 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1080_
timestamp 1649977179
transform 1 0 28520 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp 1649977179
transform 1 0 28612 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1082_
timestamp 1649977179
transform 1 0 30544 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1083_
timestamp 1649977179
transform 1 0 28612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1084_
timestamp 1649977179
transform 1 0 28336 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1085_
timestamp 1649977179
transform 1 0 25852 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1086_
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1087_
timestamp 1649977179
transform 1 0 26036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1088_
timestamp 1649977179
transform 1 0 25944 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1089_
timestamp 1649977179
transform 1 0 25668 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1090_
timestamp 1649977179
transform 1 0 23000 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1091_
timestamp 1649977179
transform 1 0 25576 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1092_
timestamp 1649977179
transform 1 0 24564 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1093_
timestamp 1649977179
transform 1 0 26036 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1094_
timestamp 1649977179
transform 1 0 25116 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1095_
timestamp 1649977179
transform 1 0 22264 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1096_
timestamp 1649977179
transform 1 0 25576 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1097_
timestamp 1649977179
transform 1 0 24932 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1098_
timestamp 1649977179
transform 1 0 22632 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1099_
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1100_
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1101_
timestamp 1649977179
transform 1 0 22632 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1102_
timestamp 1649977179
transform 1 0 23276 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1103_
timestamp 1649977179
transform 1 0 21988 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 1649977179
transform 1 0 21804 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1649977179
transform 1 0 22448 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1649977179
transform 1 0 23276 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_1  _1107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22908 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1108_
timestamp 1649977179
transform 1 0 35512 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1649977179
transform 1 0 36340 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1649977179
transform 1 0 29348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1112_
timestamp 1649977179
transform 1 0 36432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1113_
timestamp 1649977179
transform 1 0 35512 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1114_
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1115_
timestamp 1649977179
transform 1 0 36432 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1116_
timestamp 1649977179
transform 1 0 35972 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1649977179
transform 1 0 35604 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1649977179
transform 1 0 33856 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1119_
timestamp 1649977179
transform 1 0 36432 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1120_
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1121_
timestamp 1649977179
transform 1 0 33764 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1649977179
transform 1 0 33028 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1123_
timestamp 1649977179
transform 1 0 35328 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1124_
timestamp 1649977179
transform 1 0 35788 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1649977179
transform 1 0 35420 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1127_
timestamp 1649977179
transform 1 0 33396 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1128_
timestamp 1649977179
transform 1 0 35052 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1129_
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1649977179
transform 1 0 34960 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1132_
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1134_
timestamp 1649977179
transform 1 0 34776 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1135_
timestamp 1649977179
transform 1 0 34040 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1136_
timestamp 1649977179
transform 1 0 31096 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1138_
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1139_
timestamp 1649977179
transform 1 0 32108 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1140_
timestamp 1649977179
transform 1 0 31924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1141_
timestamp 1649977179
transform 1 0 33120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1142_
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1143_
timestamp 1649977179
transform 1 0 31280 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1144_
timestamp 1649977179
transform 1 0 32108 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1145_
timestamp 1649977179
transform 1 0 40112 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1146_
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1147_
timestamp 1649977179
transform 1 0 33028 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1148_
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1149_
timestamp 1649977179
transform 1 0 35604 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1150_
timestamp 1649977179
transform 1 0 36340 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1151_
timestamp 1649977179
transform 1 0 35512 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1152_
timestamp 1649977179
transform 1 0 36616 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1153_
timestamp 1649977179
transform 1 0 36064 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1154_
timestamp 1649977179
transform 1 0 36800 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1155_
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1156_
timestamp 1649977179
transform 1 0 36156 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1157_
timestamp 1649977179
transform 1 0 30728 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32384 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1159_
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1160_
timestamp 1649977179
transform 1 0 35880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1161_
timestamp 1649977179
transform 1 0 40112 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1162_
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1163_
timestamp 1649977179
transform 1 0 40756 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1164_
timestamp 1649977179
transform 1 0 37536 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1165_
timestamp 1649977179
transform 1 0 36156 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1166_
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1649977179
transform 1 0 38456 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1169_
timestamp 1649977179
transform 1 0 39192 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1170_
timestamp 1649977179
transform 1 0 38732 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1171_
timestamp 1649977179
transform 1 0 38824 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1172_
timestamp 1649977179
transform 1 0 38916 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1173_
timestamp 1649977179
transform 1 0 39652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1174_
timestamp 1649977179
transform 1 0 23828 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1649977179
transform 1 0 24656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1176_
timestamp 1649977179
transform 1 0 41124 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1649977179
transform 1 0 41216 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1178_
timestamp 1649977179
transform 1 0 41952 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1649977179
transform 1 0 42136 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1649977179
transform 1 0 42964 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1649977179
transform 1 0 44160 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1182_
timestamp 1649977179
transform 1 0 43332 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1183_
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1184_
timestamp 1649977179
transform 1 0 43792 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1185_
timestamp 1649977179
transform 1 0 46828 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1186_
timestamp 1649977179
transform 1 0 47656 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1187_
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1649977179
transform 1 0 45632 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1191_
timestamp 1649977179
transform 1 0 37352 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1192_
timestamp 1649977179
transform 1 0 38180 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 46460 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1194_
timestamp 1649977179
transform 1 0 43608 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42872 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1649977179
transform 1 0 45816 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1197_
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43792 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1199_
timestamp 1649977179
transform 1 0 45080 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1200_
timestamp 1649977179
transform 1 0 45816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1201_
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1202_
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1649977179
transform 1 0 43792 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1204_
timestamp 1649977179
transform 1 0 42780 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1205_
timestamp 1649977179
transform 1 0 43792 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1206_
timestamp 1649977179
transform 1 0 43884 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1207_
timestamp 1649977179
transform 1 0 43884 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1208_
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1649977179
transform 1 0 46736 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1210_
timestamp 1649977179
transform 1 0 45908 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1214_
timestamp 1649977179
transform 1 0 46460 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1215_
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1216_
timestamp 1649977179
transform 1 0 45724 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1217_
timestamp 1649977179
transform 1 0 44712 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1649977179
transform 1 0 45448 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 1649977179
transform 1 0 46368 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1220_
timestamp 1649977179
transform 1 0 44528 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43424 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1222_
timestamp 1649977179
transform 1 0 23092 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1649977179
transform 1 0 23644 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1649977179
transform 1 0 26128 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1225_
timestamp 1649977179
transform 1 0 24564 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1226_
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1227_
timestamp 1649977179
transform 1 0 25300 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1228_
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1229_
timestamp 1649977179
transform 1 0 24472 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1230_
timestamp 1649977179
transform 1 0 25944 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1231_
timestamp 1649977179
transform 1 0 24840 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1232_
timestamp 1649977179
transform 1 0 24196 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1233_
timestamp 1649977179
transform 1 0 24840 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1234_
timestamp 1649977179
transform 1 0 24748 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1235_
timestamp 1649977179
transform 1 0 28612 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1236_
timestamp 1649977179
transform 1 0 25760 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1237_
timestamp 1649977179
transform 1 0 25576 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1238_
timestamp 1649977179
transform 1 0 26772 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1239_
timestamp 1649977179
transform 1 0 27600 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1240_
timestamp 1649977179
transform 1 0 26772 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1241_
timestamp 1649977179
transform 1 0 25852 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1242_
timestamp 1649977179
transform 1 0 25668 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1243_
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1244_
timestamp 1649977179
transform 1 0 27048 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1245_
timestamp 1649977179
transform 1 0 27508 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1246_
timestamp 1649977179
transform 1 0 26956 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1247_
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1248_
timestamp 1649977179
transform 1 0 25944 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1250_
timestamp 1649977179
transform 1 0 26220 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1251_
timestamp 1649977179
transform 1 0 25300 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1252_
timestamp 1649977179
transform 1 0 26864 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1649977179
transform 1 0 28980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1254_
timestamp 1649977179
transform 1 0 29992 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1649977179
transform 1 0 28612 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1649977179
transform 1 0 29348 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1257_
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1649977179
transform 1 0 31464 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1260_
timestamp 1649977179
transform 1 0 32660 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1261_
timestamp 1649977179
transform 1 0 29808 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1649977179
transform 1 0 29624 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1263_
timestamp 1649977179
transform 1 0 29808 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1264_
timestamp 1649977179
transform 1 0 27600 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1265_
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1266_
timestamp 1649977179
transform 1 0 31004 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1649977179
transform 1 0 28520 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1268_
timestamp 1649977179
transform 1 0 28336 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1269_
timestamp 1649977179
transform 1 0 27968 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1270_
timestamp 1649977179
transform 1 0 28336 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1271_
timestamp 1649977179
transform 1 0 30820 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1272_
timestamp 1649977179
transform 1 0 31188 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1649977179
transform 1 0 36340 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1274_
timestamp 1649977179
transform 1 0 33212 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1649977179
transform 1 0 32476 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1276_
timestamp 1649977179
transform 1 0 33396 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1277_
timestamp 1649977179
transform 1 0 33488 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1278_
timestamp 1649977179
transform 1 0 34960 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1649977179
transform 1 0 35788 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1280_
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1649977179
transform 1 0 36432 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1282_
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1649977179
transform 1 0 37352 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1649977179
transform 1 0 38824 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1285_
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1286_
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1287_
timestamp 1649977179
transform 1 0 36984 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1288_
timestamp 1649977179
transform 1 0 34224 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1289_
timestamp 1649977179
transform 1 0 35236 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1290_
timestamp 1649977179
transform 1 0 36248 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1649977179
transform 1 0 34960 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1292_
timestamp 1649977179
transform 1 0 34776 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1293_
timestamp 1649977179
transform 1 0 40664 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1649977179
transform 1 0 40664 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 1649977179
transform 1 0 41492 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1296_
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1297_
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1649977179
transform 1 0 43240 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1299_
timestamp 1649977179
transform 1 0 43792 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1300_
timestamp 1649977179
transform 1 0 43884 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1649977179
transform 1 0 42964 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1649977179
transform 1 0 42780 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1303_
timestamp 1649977179
transform 1 0 41400 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1304_
timestamp 1649977179
transform 1 0 40020 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1305_
timestamp 1649977179
transform 1 0 40664 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1306_
timestamp 1649977179
transform 1 0 41216 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1307_
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1308_
timestamp 1649977179
transform 1 0 41492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1309_
timestamp 1649977179
transform 1 0 40756 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1310_
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1312_
timestamp 1649977179
transform 1 0 41860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1313_
timestamp 1649977179
transform 1 0 41676 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1314_
timestamp 1649977179
transform 1 0 38916 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1649977179
transform 1 0 33028 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1649977179
transform 1 0 33764 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1649977179
transform 1 0 40480 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1649977179
transform 1 0 37996 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1649977179
transform 1 0 35512 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1649977179
transform 1 0 29900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1649977179
transform 1 0 29532 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1649977179
transform 1 0 29900 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1649977179
transform 1 0 27600 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1649977179
transform 1 0 26680 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1649977179
transform 1 0 24840 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1649977179
transform 1 0 33028 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1649977179
transform 1 0 32476 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1649977179
transform 1 0 32292 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1649977179
transform 1 0 34132 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1649977179
transform 1 0 36432 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1336_
timestamp 1649977179
transform 1 0 37996 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1337_
timestamp 1649977179
transform 1 0 41400 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1649977179
transform 1 0 39836 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1649977179
transform 1 0 43148 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1340_
timestamp 1649977179
transform 1 0 36064 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1649977179
transform 1 0 46644 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1649977179
transform 1 0 46736 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1343_
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1649977179
transform 1 0 45632 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1649977179
transform 1 0 40204 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1649977179
transform 1 0 27600 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1649977179
transform 1 0 43792 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1350_
timestamp 1649977179
transform 1 0 30820 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1351_
timestamp 1649977179
transform 1 0 30912 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1352_
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1353_
timestamp 1649977179
transform 1 0 30728 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1354_
timestamp 1649977179
transform 1 0 25576 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1355_
timestamp 1649977179
transform 1 0 24840 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1356_
timestamp 1649977179
transform 1 0 23828 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1357_
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1358_
timestamp 1649977179
transform 1 0 33672 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1649977179
transform 1 0 29716 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1649977179
transform 1 0 33488 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1649977179
transform 1 0 32844 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1649977179
transform 1 0 32108 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1649977179
transform 1 0 30912 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1649977179
transform 1 0 36156 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1649977179
transform 1 0 36616 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1649977179
transform 1 0 38732 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1649977179
transform 1 0 25024 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1649977179
transform 1 0 40480 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1649977179
transform 1 0 43792 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1649977179
transform 1 0 46736 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1649977179
transform 1 0 46736 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1649977179
transform 1 0 45632 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1649977179
transform 1 0 37168 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1649977179
transform 1 0 43884 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1649977179
transform 1 0 44988 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1649977179
transform 1 0 43976 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1649977179
transform 1 0 42688 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1649977179
transform 1 0 43056 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1649977179
transform 1 0 45172 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1649977179
transform 1 0 45632 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1649977179
transform 1 0 46736 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1649977179
transform 1 0 46736 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1649977179
transform 1 0 42780 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1649977179
transform 1 0 24380 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1649977179
transform 1 0 24656 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1649977179
transform 1 0 24104 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1649977179
transform 1 0 25024 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1649977179
transform 1 0 27876 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1649977179
transform 1 0 26496 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1649977179
transform 1 0 24472 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1649977179
transform 1 0 25024 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1649977179
transform 1 0 27140 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1649977179
transform 1 0 30820 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1649977179
transform 1 0 28796 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1649977179
transform 1 0 31372 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1649977179
transform 1 0 32384 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1649977179
transform 1 0 33120 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1649977179
transform 1 0 35236 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1649977179
transform 1 0 37076 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1649977179
transform 1 0 37996 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1649977179
transform 1 0 39836 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1649977179
transform 1 0 40204 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1649977179
transform 1 0 41124 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1649977179
transform 1 0 42964 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1649977179
transform 1 0 43976 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1649977179
transform 1 0 39560 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1649977179
transform 1 0 40848 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1649977179
transform 1 0 40020 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1527__10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1528__11
timestamp 1649977179
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1649977179
transform 1 0 2116 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1529__12
timestamp 1649977179
transform 1 0 19688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1530__13
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1649977179
transform 1 0 19504 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1531__14
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1532__15
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1649977179
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1533__16
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1534__17
timestamp 1649977179
transform 1 0 4232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1535__18
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1649977179
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1649977179
transform 1 0 46276 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1536__19
timestamp 1649977179
transform 1 0 45816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1537__20
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1649977179
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1538__21
timestamp 1649977179
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1649977179
transform 1 0 21988 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1539__22
timestamp 1649977179
transform 1 0 46828 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1649977179
transform 1 0 45172 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1540__23
timestamp 1649977179
transform 1 0 4048 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1649977179
transform 1 0 3956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1541__24
timestamp 1649977179
transform 1 0 26220 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1542__25
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1543__26
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1649977179
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1649977179
transform 1 0 46276 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1544__27
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1545__28
timestamp 1649977179
transform 1 0 5336 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1545_
timestamp 1649977179
transform 1 0 5244 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1546__29
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1546_
timestamp 1649977179
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1547_
timestamp 1649977179
transform 1 0 2760 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1547__30
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1548__31
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1548_
timestamp 1649977179
transform 1 0 45172 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1549__32
timestamp 1649977179
transform 1 0 29900 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1549_
timestamp 1649977179
transform 1 0 29716 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1550_
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1550__33
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1551_
timestamp 1649977179
transform 1 0 46276 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1551__34
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1552_
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1552__35
timestamp 1649977179
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1553__36
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1553_
timestamp 1649977179
transform 1 0 46276 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1554__37
timestamp 1649977179
transform 1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1554_
timestamp 1649977179
transform 1 0 2024 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1555__38
timestamp 1649977179
transform 1 0 45632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1555_
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1556__39
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1556_
timestamp 1649977179
transform 1 0 6072 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1557__40
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1557_
timestamp 1649977179
transform 1 0 46276 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1558__41
timestamp 1649977179
transform 1 0 46184 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1558_
timestamp 1649977179
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1559__42
timestamp 1649977179
transform 1 0 27048 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1559_
timestamp 1649977179
transform 1 0 26956 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1560__43
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1560_
timestamp 1649977179
transform 1 0 32752 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1561__44
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1561_
timestamp 1649977179
transform 1 0 7728 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1562__45
timestamp 1649977179
transform 1 0 2116 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1562_
timestamp 1649977179
transform 1 0 2116 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1563__46
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1563_
timestamp 1649977179
transform 1 0 46276 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1564_
timestamp 1649977179
transform 1 0 22264 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1564__47
timestamp 1649977179
transform 1 0 22816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1565__48
timestamp 1649977179
transform 1 0 45632 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1565_
timestamp 1649977179
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1566__49
timestamp 1649977179
transform 1 0 2944 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1566_
timestamp 1649977179
transform 1 0 2116 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1567__50
timestamp 1649977179
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1567_
timestamp 1649977179
transform 1 0 18676 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1568__51
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1568_
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1569_
timestamp 1649977179
transform 1 0 46276 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1569__52
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1570_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1570__53
timestamp 1649977179
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1571__54
timestamp 1649977179
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1571_
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1572_
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1572__55
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1573_
timestamp 1649977179
transform 1 0 41492 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1574_
timestamp 1649977179
transform 1 0 21988 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1575_
timestamp 1649977179
transform 1 0 41216 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1576_
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1577__56
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1577_
timestamp 1649977179
transform 1 0 45172 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1578__57
timestamp 1649977179
transform 1 0 2116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1578_
timestamp 1649977179
transform 1 0 2024 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1579__58
timestamp 1649977179
transform 1 0 40204 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1579_
timestamp 1649977179
transform 1 0 40020 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1580_
timestamp 1649977179
transform 1 0 8832 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1580__59
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1581__60
timestamp 1649977179
transform 1 0 31556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1581_
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1582__61
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1582_
timestamp 1649977179
transform 1 0 46276 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1583__62
timestamp 1649977179
transform 1 0 27600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1583_
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1584__63
timestamp 1649977179
transform 1 0 35880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1584_
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1585__64
timestamp 1649977179
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1585_
timestamp 1649977179
transform 1 0 2392 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1586__65
timestamp 1649977179
transform 1 0 38088 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1586_
timestamp 1649977179
transform 1 0 38088 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1587__66
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1587_
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1588_
timestamp 1649977179
transform 1 0 46276 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1588__67
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1589__68
timestamp 1649977179
transform 1 0 1472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1589_
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1590__69
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1590_
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1591_
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1591__70
timestamp 1649977179
transform 1 0 1748 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1592_
timestamp 1649977179
transform 1 0 46276 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1592__71
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1593__72
timestamp 1649977179
transform 1 0 45632 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1593_
timestamp 1649977179
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1594__73
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1594_
timestamp 1649977179
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1595__74
timestamp 1649977179
transform 1 0 15456 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1595_
timestamp 1649977179
transform 1 0 15364 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1596__75
timestamp 1649977179
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1596_
timestamp 1649977179
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1597_
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1597__76
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1598__77
timestamp 1649977179
transform 1 0 39284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1598_
timestamp 1649977179
transform 1 0 38548 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1599__78
timestamp 1649977179
transform 1 0 41584 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1599_
timestamp 1649977179
transform 1 0 41584 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1600_
timestamp 1649977179
transform 1 0 25300 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1600__79
timestamp 1649977179
transform 1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1601__80
timestamp 1649977179
transform 1 0 44160 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1601_
timestamp 1649977179
transform 1 0 44712 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1602__81
timestamp 1649977179
transform 1 0 2116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1602_
timestamp 1649977179
transform 1 0 2116 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1603_
timestamp 1649977179
transform 1 0 13432 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1603__82
timestamp 1649977179
transform 1 0 12788 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1604__83
timestamp 1649977179
transform 1 0 12512 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1604_
timestamp 1649977179
transform 1 0 11868 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1605__84
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1605_
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1606__85
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1606_
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1607__86
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1607_
timestamp 1649977179
transform 1 0 2116 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1608_
timestamp 1649977179
transform 1 0 46276 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1608__87
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1609__88
timestamp 1649977179
transform 1 0 47472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1609_
timestamp 1649977179
transform 1 0 46276 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1610__89
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1610_
timestamp 1649977179
transform 1 0 46276 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1611__90
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1611_
timestamp 1649977179
transform 1 0 2116 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1612__91
timestamp 1649977179
transform 1 0 13248 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1612_
timestamp 1649977179
transform 1 0 13156 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1613__92
timestamp 1649977179
transform 1 0 44528 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1613_
timestamp 1649977179
transform 1 0 45172 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1614__93
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1614_
timestamp 1649977179
transform 1 0 13432 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1615__94
timestamp 1649977179
transform 1 0 36432 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1615_
timestamp 1649977179
transform 1 0 35696 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1616__95
timestamp 1649977179
transform 1 0 14260 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1616_
timestamp 1649977179
transform 1 0 14168 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1617_
timestamp 1649977179
transform 1 0 46276 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1617__96
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1618_
timestamp 1649977179
transform 1 0 1656 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1618__97
timestamp 1649977179
transform 1 0 2392 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1619__98
timestamp 1649977179
transform 1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1619_
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1620__99
timestamp 1649977179
transform 1 0 24656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1620_
timestamp 1649977179
transform 1 0 24656 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1621__100
timestamp 1649977179
transform 1 0 25300 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1621_
timestamp 1649977179
transform 1 0 24564 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1622_
timestamp 1649977179
transform 1 0 46276 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1622__101
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1623__102
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1623_
timestamp 1649977179
transform 1 0 46276 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1624__103
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1624_
timestamp 1649977179
transform 1 0 28612 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1625__104
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1625_
timestamp 1649977179
transform 1 0 42136 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1626__105
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1626_
timestamp 1649977179
transform 1 0 46276 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1627__106
timestamp 1649977179
transform 1 0 4692 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1627_
timestamp 1649977179
transform 1 0 2300 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1628_
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1628__107
timestamp 1649977179
transform 1 0 40848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1629__108
timestamp 1649977179
transform 1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1629_
timestamp 1649977179
transform 1 0 2116 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1630__109
timestamp 1649977179
transform 1 0 42136 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1630_
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1631__110
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1631_
timestamp 1649977179
transform 1 0 10856 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1632__111
timestamp 1649977179
transform 1 0 2116 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1632_
timestamp 1649977179
transform 1 0 2024 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1633__112
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1633_
timestamp 1649977179
transform 1 0 2024 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1634__113
timestamp 1649977179
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1634_
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36340 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1649977179
transform 1 0 31188 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1649977179
transform 1 0 26036 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1649977179
transform 1 0 39008 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1649977179
transform 1 0 41584 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1649977179
transform 1 0 39008 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1649977179
transform 1 0 41584 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1649977179
transform 1 0 1564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 27784 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1649977179
transform 1 0 47840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater9
timestamp 1649977179
transform 1 0 43240 0 1 27200
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 46188 800 46428 0 FreeSans 960 0 0 0 active
port 0 nsew signal input
flabel metal2 s 15446 0 15558 800 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 27682 49200 27794 50000 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s -10 49200 102 50000 0 FreeSans 448 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal3 s 49200 42108 50000 42348 0 FreeSans 960 0 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 23818 0 23930 800 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 18666 49200 18778 50000 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal3 s 49200 44148 50000 44388 0 FreeSans 960 0 0 0 io_in[15]
port 7 nsew signal input
flabel metal3 s 49200 4028 50000 4268 0 FreeSans 960 0 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 10294 49200 10406 50000 0 FreeSans 448 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 12226 49200 12338 50000 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 43138 0 43250 800 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal3 s 0 16268 800 16508 0 FreeSans 960 0 0 0 io_in[1]
port 12 nsew signal input
flabel metal3 s 0 29188 800 29428 0 FreeSans 960 0 0 0 io_in[20]
port 13 nsew signal input
flabel metal3 s 0 18988 800 19228 0 FreeSans 960 0 0 0 io_in[21]
port 14 nsew signal input
flabel metal3 s 49200 15588 50000 15828 0 FreeSans 960 0 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 9006 49200 9118 50000 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 6430 49200 6542 50000 0 FreeSans 448 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 37342 0 37454 800 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 36698 0 36810 800 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal3 s 49200 10828 50000 11068 0 FreeSans 960 0 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 32834 0 32946 800 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 49578 49200 49690 50000 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 16090 0 16202 800 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal3 s 49200 19668 50000 19908 0 FreeSans 960 0 0 0 io_in[30]
port 24 nsew signal input
flabel metal3 s 0 44148 800 44388 0 FreeSans 960 0 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 30902 0 31014 800 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal3 s 0 25788 800 26028 0 FreeSans 960 0 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 37986 49200 38098 50000 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 43138 49200 43250 50000 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal3 s 49200 31228 50000 31468 0 FreeSans 960 0 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 44426 49200 44538 50000 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 28970 49200 29082 50000 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal3 s 49200 30548 50000 30788 0 FreeSans 960 0 0 0 io_in[4]
port 33 nsew signal input
flabel metal3 s 49200 48228 50000 48468 0 FreeSans 960 0 0 0 io_in[5]
port 34 nsew signal input
flabel metal3 s 0 30548 800 30788 0 FreeSans 960 0 0 0 io_in[6]
port 35 nsew signal input
flabel metal3 s 0 21028 800 21268 0 FreeSans 960 0 0 0 io_in[7]
port 36 nsew signal input
flabel metal3 s 49200 33268 50000 33508 0 FreeSans 960 0 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 8362 49200 8474 50000 0 FreeSans 448 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 26394 0 26506 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal bidirectional
flabel metal3 s 0 16948 800 17188 0 FreeSans 960 0 0 0 io_oeb[10]
port 40 nsew signal bidirectional
flabel metal3 s 49200 28508 50000 28748 0 FreeSans 960 0 0 0 io_oeb[11]
port 41 nsew signal bidirectional
flabel metal3 s 49200 14908 50000 15148 0 FreeSans 960 0 0 0 io_oeb[12]
port 42 nsew signal bidirectional
flabel metal3 s 49200 13548 50000 13788 0 FreeSans 960 0 0 0 io_oeb[13]
port 43 nsew signal bidirectional
flabel metal3 s 0 4708 800 4948 0 FreeSans 960 0 0 0 io_oeb[14]
port 44 nsew signal bidirectional
flabel metal2 s 14158 49200 14270 50000 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal bidirectional
flabel metal3 s 49200 1988 50000 2228 0 FreeSans 960 0 0 0 io_oeb[16]
port 46 nsew signal bidirectional
flabel metal2 s 13514 0 13626 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal bidirectional
flabel metal2 s 36054 49200 36166 50000 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal bidirectional
flabel metal2 s 14802 49200 14914 50000 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal bidirectional
flabel metal2 s 39274 0 39386 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 50 nsew signal bidirectional
flabel metal3 s 49200 21708 50000 21948 0 FreeSans 960 0 0 0 io_oeb[20]
port 51 nsew signal bidirectional
flabel metal2 s 1922 49200 2034 50000 0 FreeSans 448 90 0 0 io_oeb[21]
port 52 nsew signal bidirectional
flabel metal2 s 5142 0 5254 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal bidirectional
flabel metal2 s 25106 49200 25218 50000 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal bidirectional
flabel metal2 s 25750 49200 25862 50000 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal bidirectional
flabel metal2 s 47646 0 47758 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 56 nsew signal bidirectional
flabel metal3 s 49200 39388 50000 39628 0 FreeSans 960 0 0 0 io_oeb[26]
port 57 nsew signal bidirectional
flabel metal2 s 29614 49200 29726 50000 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal bidirectional
flabel metal2 s 41850 0 41962 800 0 FreeSans 448 90 0 0 io_oeb[28]
port 59 nsew signal bidirectional
flabel metal3 s 49200 32588 50000 32828 0 FreeSans 960 0 0 0 io_oeb[29]
port 60 nsew signal bidirectional
flabel metal2 s 41850 49200 41962 50000 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal bidirectional
flabel metal2 s 2566 49200 2678 50000 0 FreeSans 448 90 0 0 io_oeb[30]
port 62 nsew signal bidirectional
flabel metal2 s 41206 0 41318 800 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal bidirectional
flabel metal3 s 0 25108 800 25348 0 FreeSans 960 0 0 0 io_oeb[32]
port 64 nsew signal bidirectional
flabel metal2 s 48934 0 49046 800 0 FreeSans 448 90 0 0 io_oeb[33]
port 65 nsew signal bidirectional
flabel metal2 s 10938 49200 11050 50000 0 FreeSans 448 90 0 0 io_oeb[34]
port 66 nsew signal bidirectional
flabel metal3 s 0 21708 800 21948 0 FreeSans 960 0 0 0 io_oeb[35]
port 67 nsew signal bidirectional
flabel metal3 s 0 11508 800 11748 0 FreeSans 960 0 0 0 io_oeb[36]
port 68 nsew signal bidirectional
flabel metal3 s 0 18308 800 18548 0 FreeSans 960 0 0 0 io_oeb[37]
port 69 nsew signal bidirectional
flabel metal2 s 25750 0 25862 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal bidirectional
flabel metal3 s 49200 -52 50000 188 0 FreeSans 960 0 0 0 io_oeb[4]
port 71 nsew signal bidirectional
flabel metal3 s 0 32588 800 32828 0 FreeSans 960 0 0 0 io_oeb[5]
port 72 nsew signal bidirectional
flabel metal3 s 49200 17628 50000 17868 0 FreeSans 960 0 0 0 io_oeb[6]
port 73 nsew signal bidirectional
flabel metal2 s 12870 49200 12982 50000 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal bidirectional
flabel metal2 s 4498 0 4610 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal bidirectional
flabel metal2 s 10938 0 11050 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal bidirectional
flabel metal3 s 49200 46868 50000 47108 0 FreeSans 960 0 0 0 io_out[0]
port 77 nsew signal bidirectional
flabel metal3 s 49200 27828 50000 28068 0 FreeSans 960 0 0 0 io_out[10]
port 78 nsew signal bidirectional
flabel metal3 s 0 2668 800 2908 0 FreeSans 960 0 0 0 io_out[11]
port 79 nsew signal bidirectional
flabel metal3 s 0 7428 800 7668 0 FreeSans 960 0 0 0 io_out[12]
port 80 nsew signal bidirectional
flabel metal2 s 40562 0 40674 800 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal bidirectional
flabel metal3 s 49200 40068 50000 40308 0 FreeSans 960 0 0 0 io_out[14]
port 82 nsew signal bidirectional
flabel metal3 s 0 41428 800 41668 0 FreeSans 960 0 0 0 io_out[15]
port 83 nsew signal bidirectional
flabel metal3 s 49200 26468 50000 26708 0 FreeSans 960 0 0 0 io_out[16]
port 84 nsew signal bidirectional
flabel metal2 s 46358 49200 46470 50000 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal bidirectional
flabel metal2 s 47002 0 47114 800 0 FreeSans 448 90 0 0 io_out[18]
port 86 nsew signal bidirectional
flabel metal3 s 0 23748 800 23988 0 FreeSans 960 0 0 0 io_out[19]
port 87 nsew signal bidirectional
flabel metal2 s 33478 49200 33590 50000 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal bidirectional
flabel metal2 s 40562 49200 40674 50000 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal bidirectional
flabel metal3 s 0 40748 800 40988 0 FreeSans 960 0 0 0 io_out[21]
port 90 nsew signal bidirectional
flabel metal2 s 32190 0 32302 800 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal bidirectional
flabel metal3 s 49200 22388 50000 22628 0 FreeSans 960 0 0 0 io_out[23]
port 92 nsew signal bidirectional
flabel metal2 s 27682 0 27794 800 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal bidirectional
flabel metal2 s 36698 49200 36810 50000 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal bidirectional
flabel metal3 s 0 5388 800 5628 0 FreeSans 960 0 0 0 io_out[26]
port 95 nsew signal bidirectional
flabel metal2 s 38630 49200 38742 50000 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal bidirectional
flabel metal2 s 17378 0 17490 800 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal bidirectional
flabel metal3 s 49200 1308 50000 1548 0 FreeSans 960 0 0 0 io_out[29]
port 98 nsew signal bidirectional
flabel metal2 s 7074 0 7186 800 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal bidirectional
flabel metal3 s 0 6748 800 6988 0 FreeSans 960 0 0 0 io_out[30]
port 100 nsew signal bidirectional
flabel metal3 s 0 14228 800 14468 0 FreeSans 960 0 0 0 io_out[31]
port 101 nsew signal bidirectional
flabel metal3 s 0 47548 800 47788 0 FreeSans 960 0 0 0 io_out[32]
port 102 nsew signal bidirectional
flabel metal3 s 49200 6748 50000 6988 0 FreeSans 960 0 0 0 io_out[33]
port 103 nsew signal bidirectional
flabel metal3 s 49200 41428 50000 41668 0 FreeSans 960 0 0 0 io_out[34]
port 104 nsew signal bidirectional
flabel metal3 s 49200 38028 50000 38268 0 FreeSans 960 0 0 0 io_out[35]
port 105 nsew signal bidirectional
flabel metal2 s 15446 49200 15558 50000 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal bidirectional
flabel metal3 s 49200 44828 50000 45068 0 FreeSans 960 0 0 0 io_out[37]
port 107 nsew signal bidirectional
flabel metal3 s 0 43468 800 43708 0 FreeSans 960 0 0 0 io_out[3]
port 108 nsew signal bidirectional
flabel metal3 s 49200 29188 50000 29428 0 FreeSans 960 0 0 0 io_out[4]
port 109 nsew signal bidirectional
flabel metal2 s 23174 49200 23286 50000 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal bidirectional
flabel metal2 s 48290 49200 48402 50000 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal bidirectional
flabel metal3 s 0 20348 800 20588 0 FreeSans 960 0 0 0 io_out[7]
port 112 nsew signal bidirectional
flabel metal2 s 19310 0 19422 800 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal bidirectional
flabel metal3 s 0 14908 800 15148 0 FreeSans 960 0 0 0 io_out[9]
port 114 nsew signal bidirectional
flabel metal3 s 49200 8108 50000 8348 0 FreeSans 960 0 0 0 la1_data_in[0]
port 115 nsew signal input
flabel metal2 s 21886 0 21998 800 0 FreeSans 448 90 0 0 la1_data_in[10]
port 116 nsew signal input
flabel metal3 s 49200 6068 50000 6308 0 FreeSans 960 0 0 0 la1_data_in[11]
port 117 nsew signal input
flabel metal3 s 0 37348 800 37588 0 FreeSans 960 0 0 0 la1_data_in[12]
port 118 nsew signal input
flabel metal2 s 34122 0 34234 800 0 FreeSans 448 90 0 0 la1_data_in[13]
port 119 nsew signal input
flabel metal3 s 0 13548 800 13788 0 FreeSans 960 0 0 0 la1_data_in[14]
port 120 nsew signal input
flabel metal2 s 16734 49200 16846 50000 0 FreeSans 448 90 0 0 la1_data_in[15]
port 121 nsew signal input
flabel metal2 s 31546 49200 31658 50000 0 FreeSans 448 90 0 0 la1_data_in[16]
port 122 nsew signal input
flabel metal2 s 23818 49200 23930 50000 0 FreeSans 448 90 0 0 la1_data_in[17]
port 123 nsew signal input
flabel metal2 s 43782 0 43894 800 0 FreeSans 448 90 0 0 la1_data_in[18]
port 124 nsew signal input
flabel metal2 s 17378 49200 17490 50000 0 FreeSans 448 90 0 0 la1_data_in[19]
port 125 nsew signal input
flabel metal2 s 19954 0 20066 800 0 FreeSans 448 90 0 0 la1_data_in[1]
port 126 nsew signal input
flabel metal3 s 0 36668 800 36908 0 FreeSans 960 0 0 0 la1_data_in[20]
port 127 nsew signal input
flabel metal2 s 48934 49200 49046 50000 0 FreeSans 448 90 0 0 la1_data_in[21]
port 128 nsew signal input
flabel metal3 s 49200 8788 50000 9028 0 FreeSans 960 0 0 0 la1_data_in[22]
port 129 nsew signal input
flabel metal3 s 0 628 800 868 0 FreeSans 960 0 0 0 la1_data_in[23]
port 130 nsew signal input
flabel metal2 s 14158 0 14270 800 0 FreeSans 448 90 0 0 la1_data_in[24]
port 131 nsew signal input
flabel metal3 s 0 38708 800 38948 0 FreeSans 960 0 0 0 la1_data_in[25]
port 132 nsew signal input
flabel metal3 s 49200 3348 50000 3588 0 FreeSans 960 0 0 0 la1_data_in[26]
port 133 nsew signal input
flabel metal2 s 28970 0 29082 800 0 FreeSans 448 90 0 0 la1_data_in[27]
port 134 nsew signal input
flabel metal3 s 0 33948 800 34188 0 FreeSans 960 0 0 0 la1_data_in[28]
port 135 nsew signal input
flabel metal2 s 1278 49200 1390 50000 0 FreeSans 448 90 0 0 la1_data_in[29]
port 136 nsew signal input
flabel metal2 s 11582 0 11694 800 0 FreeSans 448 90 0 0 la1_data_in[2]
port 137 nsew signal input
flabel metal2 s 1278 0 1390 800 0 FreeSans 448 90 0 0 la1_data_in[30]
port 138 nsew signal input
flabel metal2 s 38630 0 38742 800 0 FreeSans 448 90 0 0 la1_data_in[31]
port 139 nsew signal input
flabel metal3 s 0 31908 800 32148 0 FreeSans 960 0 0 0 la1_data_in[3]
port 140 nsew signal input
flabel metal2 s 42494 49200 42606 50000 0 FreeSans 448 90 0 0 la1_data_in[4]
port 141 nsew signal input
flabel metal3 s 49200 24428 50000 24668 0 FreeSans 960 0 0 0 la1_data_in[5]
port 142 nsew signal input
flabel metal2 s 19310 49200 19422 50000 0 FreeSans 448 90 0 0 la1_data_in[6]
port 143 nsew signal input
flabel metal3 s 0 23068 800 23308 0 FreeSans 960 0 0 0 la1_data_in[7]
port 144 nsew signal input
flabel metal2 s 20598 49200 20710 50000 0 FreeSans 448 90 0 0 la1_data_in[8]
port 145 nsew signal input
flabel metal3 s 0 34628 800 34868 0 FreeSans 960 0 0 0 la1_data_in[9]
port 146 nsew signal input
flabel metal2 s 7718 0 7830 800 0 FreeSans 448 90 0 0 la1_data_out[0]
port 147 nsew signal bidirectional
flabel metal3 s 49200 12188 50000 12428 0 FreeSans 960 0 0 0 la1_data_out[10]
port 148 nsew signal bidirectional
flabel metal2 s 22530 0 22642 800 0 FreeSans 448 90 0 0 la1_data_out[11]
port 149 nsew signal bidirectional
flabel metal3 s 49200 46188 50000 46428 0 FreeSans 960 0 0 0 la1_data_out[12]
port 150 nsew signal bidirectional
flabel metal2 s 4498 49200 4610 50000 0 FreeSans 448 90 0 0 la1_data_out[13]
port 151 nsew signal bidirectional
flabel metal2 s 27038 49200 27150 50000 0 FreeSans 448 90 0 0 la1_data_out[14]
port 152 nsew signal bidirectional
flabel metal3 s 0 1308 800 1548 0 FreeSans 960 0 0 0 la1_data_out[15]
port 153 nsew signal bidirectional
flabel metal3 s 49200 16948 50000 17188 0 FreeSans 960 0 0 0 la1_data_out[16]
port 154 nsew signal bidirectional
flabel metal3 s 49200 35988 50000 36228 0 FreeSans 960 0 0 0 la1_data_out[17]
port 155 nsew signal bidirectional
flabel metal2 s 5786 49200 5898 50000 0 FreeSans 448 90 0 0 la1_data_out[18]
port 156 nsew signal bidirectional
flabel metal3 s 49200 25788 50000 26028 0 FreeSans 960 0 0 0 la1_data_out[19]
port 157 nsew signal bidirectional
flabel metal3 s 0 45508 800 45748 0 FreeSans 960 0 0 0 la1_data_out[1]
port 158 nsew signal bidirectional
flabel metal3 s 0 10148 800 10388 0 FreeSans 960 0 0 0 la1_data_out[20]
port 159 nsew signal bidirectional
flabel metal3 s 49200 42788 50000 43028 0 FreeSans 960 0 0 0 la1_data_out[21]
port 160 nsew signal bidirectional
flabel metal2 s 30258 49200 30370 50000 0 FreeSans 448 90 0 0 la1_data_out[22]
port 161 nsew signal bidirectional
flabel metal2 s 12870 0 12982 800 0 FreeSans 448 90 0 0 la1_data_out[23]
port 162 nsew signal bidirectional
flabel metal3 s 49200 18988 50000 19228 0 FreeSans 960 0 0 0 la1_data_out[24]
port 163 nsew signal bidirectional
flabel metal3 s 0 3348 800 3588 0 FreeSans 960 0 0 0 la1_data_out[25]
port 164 nsew signal bidirectional
flabel metal3 s 49200 5388 50000 5628 0 FreeSans 960 0 0 0 la1_data_out[26]
port 165 nsew signal bidirectional
flabel metal3 s 0 48228 800 48468 0 FreeSans 960 0 0 0 la1_data_out[27]
port 166 nsew signal bidirectional
flabel metal2 s 45070 0 45182 800 0 FreeSans 448 90 0 0 la1_data_out[28]
port 167 nsew signal bidirectional
flabel metal2 s 6430 0 6542 800 0 FreeSans 448 90 0 0 la1_data_out[29]
port 168 nsew signal bidirectional
flabel metal2 s 20598 0 20710 800 0 FreeSans 448 90 0 0 la1_data_out[2]
port 169 nsew signal bidirectional
flabel metal3 s 49200 12868 50000 13108 0 FreeSans 960 0 0 0 la1_data_out[30]
port 170 nsew signal bidirectional
flabel metal3 s 49200 48908 50000 49148 0 FreeSans 960 0 0 0 la1_data_out[31]
port 171 nsew signal bidirectional
flabel metal3 s 0 9468 800 9708 0 FreeSans 960 0 0 0 la1_data_out[3]
port 172 nsew signal bidirectional
flabel metal2 s 45714 0 45826 800 0 FreeSans 448 90 0 0 la1_data_out[4]
port 173 nsew signal bidirectional
flabel metal2 s 3210 0 3322 800 0 FreeSans 448 90 0 0 la1_data_out[5]
port 174 nsew signal bidirectional
flabel metal3 s 49200 20348 50000 20588 0 FreeSans 960 0 0 0 la1_data_out[6]
port 175 nsew signal bidirectional
flabel metal2 s 634 0 746 800 0 FreeSans 448 90 0 0 la1_data_out[7]
port 176 nsew signal bidirectional
flabel metal3 s 49200 37348 50000 37588 0 FreeSans 960 0 0 0 la1_data_out[8]
port 177 nsew signal bidirectional
flabel metal2 s 47002 49200 47114 50000 0 FreeSans 448 90 0 0 la1_data_out[9]
port 178 nsew signal bidirectional
flabel metal2 s 49578 0 49690 800 0 FreeSans 448 90 0 0 la1_oenb[0]
port 179 nsew signal input
flabel metal2 s 45070 49200 45182 50000 0 FreeSans 448 90 0 0 la1_oenb[10]
port 180 nsew signal input
flabel metal3 s 0 27828 800 28068 0 FreeSans 960 0 0 0 la1_oenb[11]
port 181 nsew signal input
flabel metal3 s 0 29868 800 30108 0 FreeSans 960 0 0 0 la1_oenb[12]
port 182 nsew signal input
flabel metal2 s 30258 0 30370 800 0 FreeSans 448 90 0 0 la1_oenb[13]
port 183 nsew signal input
flabel metal2 s -10 0 102 800 0 FreeSans 448 90 0 0 la1_oenb[14]
port 184 nsew signal input
flabel metal2 s 35410 0 35522 800 0 FreeSans 448 90 0 0 la1_oenb[15]
port 185 nsew signal input
flabel metal3 s 0 35988 800 36228 0 FreeSans 960 0 0 0 la1_oenb[16]
port 186 nsew signal input
flabel metal2 s 3854 49200 3966 50000 0 FreeSans 448 90 0 0 la1_oenb[17]
port 187 nsew signal input
flabel metal2 s 21886 49200 21998 50000 0 FreeSans 448 90 0 0 la1_oenb[18]
port 188 nsew signal input
flabel metal3 s 0 27148 800 27388 0 FreeSans 960 0 0 0 la1_oenb[19]
port 189 nsew signal input
flabel metal2 s 9006 0 9118 800 0 FreeSans 448 90 0 0 la1_oenb[1]
port 190 nsew signal input
flabel metal2 s 2566 0 2678 800 0 FreeSans 448 90 0 0 la1_oenb[20]
port 191 nsew signal input
flabel metal2 s 32190 49200 32302 50000 0 FreeSans 448 90 0 0 la1_oenb[21]
port 192 nsew signal input
flabel metal2 s 21242 49200 21354 50000 0 FreeSans 448 90 0 0 la1_oenb[22]
port 193 nsew signal input
flabel metal2 s 24462 0 24574 800 0 FreeSans 448 90 0 0 la1_oenb[23]
port 194 nsew signal input
flabel metal2 s 39918 49200 40030 50000 0 FreeSans 448 90 0 0 la1_oenb[24]
port 195 nsew signal input
flabel metal3 s 49200 10148 50000 10388 0 FreeSans 960 0 0 0 la1_oenb[25]
port 196 nsew signal input
flabel metal3 s 0 39388 800 39628 0 FreeSans 960 0 0 0 la1_oenb[26]
port 197 nsew signal input
flabel metal3 s 49200 35308 50000 35548 0 FreeSans 960 0 0 0 la1_oenb[27]
port 198 nsew signal input
flabel metal2 s 9650 0 9762 800 0 FreeSans 448 90 0 0 la1_oenb[28]
port 199 nsew signal input
flabel metal2 s 18022 0 18134 800 0 FreeSans 448 90 0 0 la1_oenb[29]
port 200 nsew signal input
flabel metal3 s 0 8108 800 8348 0 FreeSans 960 0 0 0 la1_oenb[2]
port 201 nsew signal input
flabel metal3 s 49200 34628 50000 34868 0 FreeSans 960 0 0 0 la1_oenb[30]
port 202 nsew signal input
flabel metal2 s 28326 0 28438 800 0 FreeSans 448 90 0 0 la1_oenb[31]
port 203 nsew signal input
flabel metal2 s 35410 49200 35522 50000 0 FreeSans 448 90 0 0 la1_oenb[3]
port 204 nsew signal input
flabel metal2 s 34122 49200 34234 50000 0 FreeSans 448 90 0 0 la1_oenb[4]
port 205 nsew signal input
flabel metal3 s 0 49588 800 49828 0 FreeSans 960 0 0 0 la1_oenb[5]
port 206 nsew signal input
flabel metal2 s 7718 49200 7830 50000 0 FreeSans 448 90 0 0 la1_oenb[6]
port 207 nsew signal input
flabel metal2 s 34766 0 34878 800 0 FreeSans 448 90 0 0 la1_oenb[7]
port 208 nsew signal input
flabel metal3 s 0 12188 800 12428 0 FreeSans 960 0 0 0 la1_oenb[8]
port 209 nsew signal input
flabel metal3 s 0 42788 800 43028 0 FreeSans 960 0 0 0 la1_oenb[9]
port 210 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 211 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 212 nsew ground bidirectional
flabel metal3 s 49200 23748 50000 23988 0 FreeSans 960 0 0 0 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
